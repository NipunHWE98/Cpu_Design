module divider(input[30:0]D,
								 input[30:0]d,
								 output[31:0]q);

wire[30:0]dout,sout,sin,sp;
wire[31:0]dout1,sout1,sin1,sp1,dout2,sout2,sin2,sp2,dout3,sout3,sin3,sp3,dout4,sout4,sin4,sp4,dout5,sout5,sin5,sp5,dout6,sout6,sin6,sp6,dout7,sout7,sin7,sp7,dout8,sout8,sin8,sp8, dout9,
sout9,sin9,sp9, dout10,sout10,sin10,sp10, dout11,sout11,sin11,sp11, dout12,sout12,sin12,sp12, dout13,sout13,sin13,sp13, dout14,sout14,sin14,sp14, dout15,sout15,sin15,sp15, dout16,sout16,
sin16,sp16, dout17,sout17,sin17,sp17, dout18,sout18,sin18,sp18, dout19,sout19,sin19,sp19, dout20,sout20,sin20,sp20, dout21,sout21,sin21,sp21, dout22,sout22,sin22,sp22, dout23,sout23,sin23,sp23,
 dout24,sout24,sin24,sp24, dout25,sout25,sin25,sp25, dout26,sout26,sin26,sp26, dout27,sout27,sin27,sp27, dout28,sout28,sin28,sp28, dout29,sout29,sin29,sp29, dout30,sout30,sin30,sp30, dout31,sout31,sin31,sp31, dout32,sout32,sin32,sp32;								 

//can be implemented using a 32 bit register and clock as theres no internal clock impmentede in alu 
divide_module m00(D[30],d[0],1'b0,sp[1],dout[0],sout[0],sp[0]);
divide_module m01(1'b0,d[1],dout[0],sp[2],dout[1],sout[1],sp[1]);
divide_module m02(1'b0,d[2],dout[1],sp[3],dout[2],sout[2],sp[2]);
divide_module m03(1'b0,d[3],dout[2],sp[4],dout[3],sout[3],sp[3]);
divide_module m04(1'b0,d[4],dout[3],sp[5],dout[4],sout[4],sp[4]);
divide_module m05(1'b0,d[5],dout[4],sp[6],dout[5],sout[5],sp[5]);
divide_module m06(1'b0,d[6],dout[5],sp[7],dout[6],sout[6],sp[6]);
divide_module m07(1'b0,d[7],dout[6],sp[8],dout[7],sout[7],sp[7]);
divide_module m08(1'b0,d[8],dout[7],sp[9],dout[8],sout[8],sp[8]);
divide_module m09(1'b0,d[9],dout[8],sp[10],dout[9],sout[9],sp[9]);
divide_module m10(1'b0,d[10],dout[9],sp[11],dout[10],sout[10],sp[10]);
divide_module m11(1'b0,d[11],dout[10],sp[12],dout[11],sout[11],sp[11]);
divide_module m12(1'b0,d[12],dout[11],sp[13],dout[12],sout[12],sp[12]);
divide_module m13(1'b0,d[13],dout[12],sp[14],dout[13],sout[13],sp[13]);
divide_module m14(1'b0,d[14],dout[13],sp[15],dout[14],sout[14],sp[14]);
divide_module m15(1'b0,d[15],dout[14],sp[16],dout[15],sout[15],sp[15]);
divide_module m16(1'b0,d[16],dout[15],sp[17],dout[16],sout[16],sp[16]);
divide_module m17(1'b0,d[17],dout[16],sp[18],dout[17],sout[17],sp[17]);
divide_module m18(1'b0,d[18],dout[17],sp[19],dout[18],sout[18],sp[18]);
divide_module m19(1'b0,d[19],dout[18],sp[20],dout[19],sout[19],sp[19]);
divide_module m20(1'b0,d[20],dout[19],sp[21],dout[20],sout[20],sp[20]);
divide_module m21(1'b0,d[21],dout[20],sp[22],dout[21],sout[21],sp[21]);
divide_module m22(1'b0,d[22],dout[21],sp[23],dout[22],sout[22],sp[22]);
divide_module m23(1'b0,d[23],dout[22],sp[24],dout[23],sout[23],sp[23]);
divide_module m24(1'b0,d[24],dout[23],sp[25],dout[24],sout[24],sp[24]);
divide_module m25(1'b0,d[25],dout[24],sp[26],dout[25],sout[25],sp[25]);
divide_module m26(1'b0,d[26],dout[25],sp[27],dout[26],sout[26],sp[26]);
divide_module m27(1'b0,d[27],dout[26],sp[28],dout[27],sout[27],sp[27]);
divide_module m28(1'b0,d[28],dout[27],sp[29],dout[28],sout[28],sp[28]);
divide_module m29(1'b0,d[29],dout[28],sp[30],dout[29],sout[29],sp[29]);
divide_module m30(1'b0,d[30],dout[29],~dout[30],dout[30],sout[30],sp[30]);

divide_module m40(D[29],d[0],1'b0,sp1[1],dout1[0],sout1[0],sp1[0]);
divide_module m41(1'b0,d[1],dout1[0],sp1[2],dout1[1],sout1[1],sp1[1]);
divide_module m42(1'b0,d[2],dout1[1],sp1[3],dout1[2],sout1[2],sp1[2]);
divide_module m43(1'b0,d[3],dout1[2],sp1[4],dout1[3],sout1[3],sp1[3]);
divide_module m44(1'b0,d[4],dout1[3],sp1[5],dout1[4],sout1[4],sp1[4]);
divide_module m45(1'b0,d[5],dout1[4],sp1[6],dout1[5],sout1[5],sp1[5]);
divide_module m46(1'b0,d[6],dout1[5],sp1[7],dout1[6],sout1[6],sp1[6]);
divide_module m47(1'b0,d[7],dout1[6],sp1[8],dout1[7],sout1[7],sp1[7]);
divide_module m48(1'b0,d[8],dout1[7],sp1[9],dout1[8],sout1[8],sp1[8]);
divide_module m49(1'b0,d[9],dout1[8],sp1[10],dout1[9],sout1[9],sp1[9]);
divide_module m50(1'b0,d[10],dout1[9],sp1[11],dout1[10],sout1[10],sp1[10]);
divide_module m51(1'b0,d[11],dout1[10],sp1[12],dout1[11],sout1[11],sp1[11]);
divide_module m52(1'b0,d[12],dout1[11],sp1[13],dout1[12],sout1[12],sp1[12]);
divide_module m53(1'b0,d[13],dout1[12],sp1[14],dout1[13],sout1[13],sp1[13]);
divide_module m54(1'b0,d[14],dout1[13],sp1[15],dout1[14],sout1[14],sp1[14]);
divide_module m55(1'b0,d[15],dout1[14],sp1[16],dout1[15],sout1[15],sp1[15]);
divide_module m56(1'b0,d[16],dout1[15],sp1[17],dout1[16],sout1[16],sp1[16]);
divide_module m57(1'b0,d[17],dout1[16],sp1[18],dout1[17],sout1[17],sp1[17]);
divide_module m58(1'b0,d[18],dout1[17],sp1[19],dout1[18],sout1[18],sp1[18]);
divide_module m59(1'b0,d[19],dout1[18],sp1[20],dout1[19],sout1[19],sp1[19]);
divide_module m60(1'b0,d[20],dout1[19],sp1[21],dout1[20],sout1[20],sp1[20]);
divide_module m61(1'b0,d[21],dout1[20],sp1[22],dout1[21],sout1[21],sp1[21]);
divide_module m62(1'b0,d[22],dout1[21],sp1[23],dout1[22],sout1[22],sp1[22]);
divide_module m63(1'b0,d[23],dout1[22],sp1[24],dout1[23],sout1[23],sp1[23]);
divide_module m64(1'b0,d[24],dout1[23],sp1[25],dout1[24],sout1[24],sp1[24]);
divide_module m65(1'b0,d[25],dout1[24],sp1[26],dout1[25],sout1[25],sp1[25]);
divide_module m66(1'b0,d[26],dout1[25],sp1[27],dout1[26],sout1[26],sp1[26]);
divide_module m67(1'b0,d[27],dout1[26],sp1[28],dout1[27],sout1[27],sp1[27]);
divide_module m68(1'b0,d[28],dout1[27],sp1[29],dout1[28],sout1[28],sp1[28]);
divide_module m69(1'b0,d[29],dout1[28],sp1[30],dout1[29],sout1[29],sp1[29]);
divide_module m70(1'b0,d[30],dout1[29],~dout1[30],dout1[30],sout1[30],sp1[30]);

divide_module m8000(D[28],d[0],1'b0,sp2[1],dout2[0],sout2[0],sp2[0]);
divide_module m81(1'b0,d[1],dout2[0],sp2[2],dout2[1],sout2[1],sp2[1]);
divide_module m82(1'b0,d[2],dout2[1],sp2[3],dout2[2],sout2[2],sp2[2]);
divide_module m83(1'b0,d[3],dout2[2],sp2[4],dout2[3],sout2[3],sp2[3]);
divide_module m84(1'b0,d[4],dout2[3],sp2[5],dout2[4],sout2[4],sp2[4]);
divide_module m85(1'b0,d[5],dout2[4],sp2[6],dout2[5],sout2[5],sp2[5]);
divide_module m86(1'b0,d[6],dout2[5],sp2[7],dout2[6],sout2[6],sp2[6]);
divide_module m87(1'b0,d[7],dout2[6],sp2[8],dout2[7],sout2[7],sp2[7]);
divide_module m88(1'b0,d[8],dout2[7],sp2[9],dout2[8],sout2[8],sp2[8]);
divide_module m89(1'b0,d[9],dout2[8],sp2[10],dout2[9],sout2[9],sp2[9]);
divide_module m90(1'b0,d[10],dout2[9],sp2[11],dout2[10],sout2[10],sp2[10]);
divide_module m91(1'b0,d[11],dout2[10],sp2[12],dout2[11],sout2[11],sp2[11]);
divide_module m92(1'b0,d[12],dout2[11],sp2[13],dout2[12],sout2[12],sp2[12]);
divide_module m93(1'b0,d[13],dout2[12],sp2[14],dout2[13],sout2[13],sp2[13]);
divide_module m94(1'b0,d[14],dout2[13],sp2[15],dout2[14],sout2[14],sp2[14]);
divide_module m95(1'b0,d[15],dout2[14],sp2[16],dout2[15],sout2[15],sp2[15]);
divide_module m96(1'b0,d[16],dout2[15],sp2[17],dout2[16],sout2[16],sp2[16]);
divide_module m97(1'b0,d[17],dout2[16],sp2[18],dout2[17],sout2[17],sp2[17]);
divide_module m98(1'b0,d[18],dout2[17],sp2[19],dout2[18],sout2[18],sp2[18]);
divide_module m99(1'b0,d[19],dout2[18],sp2[20],dout2[19],sout2[19],sp2[19]);
divide_module m100(1'b0,d[20],dout2[19],sp2[21],dout2[20],sout2[20],sp2[20]);
divide_module m101(1'b0,d[21],dout2[20],sp2[22],dout2[21],sout2[21],sp2[21]);
divide_module m102(1'b0,d[22],dout2[21],sp2[23],dout2[22],sout2[22],sp2[22]);
divide_module m103(1'b0,d[23],dout2[22],sp2[24],dout2[23],sout2[23],sp2[23]);
divide_module m104(1'b0,d[24],dout2[23],sp2[25],dout2[24],sout2[24],sp2[24]);
divide_module m105(1'b0,d[25],dout2[24],sp2[26],dout2[25],sout2[25],sp2[25]);
divide_module m106(1'b0,d[26],dout2[25],sp2[27],dout2[26],sout2[26],sp2[26]);
divide_module m107(1'b0,d[27],dout2[26],sp2[28],dout2[27],sout2[27],sp2[27]);
divide_module m108(1'b0,d[28],dout2[27],sp2[29],dout2[28],sout2[28],sp2[28]);
divide_module m109(1'b0,d[29],dout2[28],sp2[30],dout2[29],sout2[29],sp2[29]);
divide_module m110(1'b0,d[30],dout2[29],~dout2[30],dout2[30],sout2[30],sp2[30]);

divide_module m120(D[27],d[0],1'b0,sp3[1],dout3[0],sout3[0],sp3[0]);
divide_module m121(1'b0,d[1],dout3[0],sp3[2],dout3[1],sout3[1],sp3[1]);
divide_module m122(1'b0,d[2],dout3[1],sp3[3],dout3[2],sout3[2],sp3[2]);
divide_module m123(1'b0,d[3],dout3[2],sp3[4],dout3[3],sout3[3],sp3[3]);
divide_module m124(1'b0,d[4],dout3[3],sp3[5],dout3[4],sout3[4],sp3[4]);
divide_module m125(1'b0,d[5],dout3[4],sp3[6],dout3[5],sout3[5],sp3[5]);
divide_module m126(1'b0,d[6],dout3[5],sp3[7],dout3[6],sout3[6],sp3[6]);
divide_module m127(1'b0,d[7],dout3[6],sp3[8],dout3[7],sout3[7],sp3[7]);
divide_module m128(1'b0,d[8],dout3[7],sp3[9],dout3[8],sout3[8],sp3[8]);
divide_module m129(1'b0,d[9],dout3[8],sp3[10],dout3[9],sout3[9],sp3[9]);
divide_module m130(1'b0,d[10],dout3[9],sp3[11],dout3[10],sout3[10],sp3[10]);
divide_module m131(1'b0,d[11],dout3[10],sp3[12],dout3[11],sout3[11],sp3[11]);
divide_module m132(1'b0,d[12],dout3[11],sp3[13],dout3[12],sout3[12],sp3[12]);
divide_module m133(1'b0,d[13],dout3[12],sp3[14],dout3[13],sout3[13],sp3[13]);
divide_module m134(1'b0,d[14],dout3[13],sp3[15],dout3[14],sout3[14],sp3[14]);
divide_module m135(1'b0,d[15],dout3[14],sp3[16],dout3[15],sout3[15],sp3[15]);
divide_module m136(1'b0,d[16],dout3[15],sp3[17],dout3[16],sout3[16],sp3[16]);
divide_module m137(1'b0,d[17],dout3[16],sp3[18],dout3[17],sout3[17],sp3[17]);
divide_module m138(1'b0,d[18],dout3[17],sp3[19],dout3[18],sout3[18],sp3[18]);
divide_module m139(1'b0,d[19],dout3[18],sp3[20],dout3[19],sout3[19],sp3[19]);
divide_module m140(1'b0,d[20],dout3[19],sp3[21],dout3[20],sout3[20],sp3[20]);
divide_module m141(1'b0,d[21],dout3[20],sp3[22],dout3[21],sout3[21],sp3[21]);
divide_module m142(1'b0,d[22],dout3[21],sp3[23],dout3[22],sout3[22],sp3[22]);
divide_module m143(1'b0,d[23],dout3[22],sp3[24],dout3[23],sout3[23],sp3[23]);
divide_module m144(1'b0,d[24],dout3[23],sp3[25],dout3[24],sout3[24],sp3[24]);
divide_module m145(1'b0,d[25],dout3[24],sp3[26],dout3[25],sout3[25],sp3[25]);
divide_module m146(1'b0,d[26],dout3[25],sp3[27],dout3[26],sout3[26],sp3[26]);
divide_module m147(1'b0,d[27],dout3[26],sp3[28],dout3[27],sout3[27],sp3[27]);
divide_module m148(1'b0,d[28],dout3[27],sp3[29],dout3[28],sout3[28],sp3[28]);
divide_module m149(1'b0,d[29],dout3[28],sp3[30],dout3[29],sout3[29],sp3[29]);
divide_module m150(1'b0,d[30],dout3[29],~dout3[30],dout3[30],sout3[30],sp3[30]);


divide_module m160(D[26],d[0],1'b0,sp4[1],dout4[0],sout4[0],sp4[0]);
divide_module m161(1'b0,d[1],dout4[0],sp4[2],dout4[1],sout4[1],sp4[1]);
divide_module m162(1'b0,d[2],dout4[1],sp4[3],dout4[2],sout4[2],sp4[2]);
divide_module m163(1'b0,d[3],dout4[2],sp4[4],dout4[3],sout4[3],sp4[3]);
divide_module m164(1'b0,d[4],dout4[3],sp4[5],dout4[4],sout4[4],sp4[4]);
divide_module m165(1'b0,d[5],dout4[4],sp4[6],dout4[5],sout4[5],sp4[5]);
divide_module m166(1'b0,d[6],dout4[5],sp4[7],dout4[6],sout4[6],sp4[6]);
divide_module m167(1'b0,d[7],dout4[6],sp4[8],dout4[7],sout4[7],sp4[7]);
divide_module m168(1'b0,d[8],dout4[7],sp4[9],dout4[8],sout4[8],sp4[8]);
divide_module m169(1'b0,d[9],dout4[8],sp4[10],dout4[9],sout4[9],sp4[9]);
divide_module m170(1'b0,d[10],dout4[9],sp4[11],dout4[10],sout4[10],sp4[10]);
divide_module m171(1'b0,d[11],dout4[10],sp4[12],dout4[11],sout4[11],sp4[11]);
divide_module m172(1'b0,d[12],dout4[11],sp4[13],dout4[12],sout4[12],sp4[12]);
divide_module m173(1'b0,d[13],dout4[12],sp4[14],dout4[13],sout4[13],sp4[13]);
divide_module m174(1'b0,d[14],dout4[13],sp4[15],dout4[14],sout4[14],sp4[14]);
divide_module m175(1'b0,d[15],dout4[14],sp4[16],dout4[15],sout4[15],sp4[15]);
divide_module m176(1'b0,d[16],dout4[15],sp4[17],dout4[16],sout4[16],sp4[16]);
divide_module m177(1'b0,d[17],dout4[16],sp4[18],dout4[17],sout4[17],sp4[17]);
divide_module m178(1'b0,d[18],dout4[17],sp4[19],dout4[18],sout4[18],sp4[18]);
divide_module m179(1'b0,d[19],dout4[18],sp4[20],dout4[19],sout4[19],sp4[19]);
divide_module m180(1'b0,d[20],dout4[19],sp4[21],dout4[20],sout4[20],sp4[20]);
divide_module m181(1'b0,d[21],dout4[20],sp4[22],dout4[21],sout4[21],sp4[21]);
divide_module m182(1'b0,d[22],dout4[21],sp4[23],dout4[22],sout4[22],sp4[22]);
divide_module m183(1'b0,d[23],dout4[22],sp4[24],dout4[23],sout4[23],sp4[23]);
divide_module m184(1'b0,d[24],dout4[23],sp4[25],dout4[24],sout4[24],sp4[24]);
divide_module m185(1'b0,d[25],dout4[24],sp4[26],dout4[25],sout4[25],sp4[25]);
divide_module m186(1'b0,d[26],dout4[25],sp4[27],dout4[26],sout4[26],sp4[26]);
divide_module m187(1'b0,d[27],dout4[26],sp4[28],dout4[27],sout4[27],sp4[27]);
divide_module m188(1'b0,d[28],dout4[27],sp4[29],dout4[28],sout4[28],sp4[28]);
divide_module m189(1'b0,d[29],dout4[28],sp4[30],dout4[29],sout4[29],sp4[29]);
divide_module m190(1'b0,d[30],dout4[29],~dout4[30],dout4[30],sout4[30],sp4[30]);

divide_module m1600(D[25],d[0],1'b0,sp5[1],dout5[0],sout5[0],sp5[0]);
divide_module m1610(1'b0,d[1],dout5[0],sp5[2],dout5[1],sout5[1],sp5[1]);
divide_module m1620(1'b0,d[2],dout5[1],sp5[3],dout5[2],sout5[2],sp5[2]);
divide_module m1630(1'b0,d[3],dout5[2],sp5[4],dout5[3],sout5[3],sp5[3]);
divide_module m1640(1'b0,d[4],dout5[3],sp5[5],dout5[4],sout5[4],sp5[4]);
divide_module m1650(1'b0,d[5],dout5[4],sp5[6],dout5[5],sout5[5],sp5[5]);
divide_module m1660(1'b0,d[6],dout5[5],sp5[7],dout5[6],sout5[6],sp5[6]);
divide_module m1670(1'b0,d[7],dout5[6],sp5[8],dout5[7],sout5[7],sp5[7]);
divide_module m1680(1'b0,d[8],dout5[7],sp5[9],dout5[8],sout5[8],sp5[8]);
divide_module m1690(1'b0,d[9],dout5[8],sp5[10],dout5[9],sout5[9],sp5[9]);
divide_module m1700(1'b0,d[10],dout5[9],sp5[11],dout5[10],sout5[10],sp5[10]);
divide_module m1710(1'b0,d[11],dout5[10],sp5[12],dout5[11],sout5[11],sp5[11]);
divide_module m1720(1'b0,d[12],dout5[11],sp5[13],dout5[12],sout5[12],sp5[12]);
divide_module m1730(1'b0,d[13],dout5[12],sp5[14],dout5[13],sout5[13],sp5[13]);
divide_module m1740(1'b0,d[14],dout5[13],sp5[15],dout5[14],sout5[14],sp5[14]);
divide_module m1750(1'b0,d[15],dout5[14],sp5[16],dout5[15],sout5[15],sp5[15]);
divide_module m1760(1'b0,d[16],dout5[15],sp5[17],dout5[16],sout5[16],sp5[16]);
divide_module m1770(1'b0,d[17],dout5[16],sp5[18],dout5[17],sout5[17],sp5[17]);
divide_module m1780(1'b0,d[18],dout5[17],sp5[19],dout5[18],sout5[18],sp5[18]);
divide_module m1790(1'b0,d[19],dout5[18],sp5[20],dout5[19],sout5[19],sp5[19]);
divide_module m1800(1'b0,d[20],dout5[19],sp5[21],dout5[20],sout5[20],sp5[20]);
divide_module m1810(1'b0,d[21],dout5[20],sp5[22],dout5[21],sout5[21],sp5[21]);
divide_module m1820(1'b0,d[22],dout5[21],sp5[23],dout5[22],sout5[22],sp5[22]);
divide_module m1830(1'b0,d[23],dout5[22],sp5[24],dout5[23],sout5[23],sp5[23]);
divide_module m1840(1'b0,d[24],dout5[23],sp5[25],dout5[24],sout5[24],sp5[24]);
divide_module m1850(1'b0,d[25],dout5[24],sp5[26],dout5[25],sout5[25],sp5[25]);
divide_module m1860(1'b0,d[26],dout5[25],sp5[27],dout5[26],sout5[26],sp5[26]);
divide_module m1870(1'b0,d[27],dout5[26],sp5[28],dout5[27],sout5[27],sp5[27]);
divide_module m1880(1'b0,d[28],dout5[27],sp5[29],dout5[28],sout5[28],sp5[28]);
divide_module m1890(1'b0,d[29],dout5[28],sp5[30],dout5[29],sout5[29],sp5[29]);
divide_module m1900(1'b0,d[30],dout5[29],~dout5[30],dout5[30],sout5[30],sp5[30]);

divide_module m1601(D[24],d[0],1'b0,sp6[1],dout6[0],sout6[0],sp6[0]);
divide_module m1611(1'b0,d[1],dout6[0],sp6[2],dout6[1],sout6[1],sp6[1]);
divide_module m1621(1'b0,d[2],dout6[1],sp6[3],dout6[2],sout6[2],sp6[2]);
divide_module m1631(1'b0,d[3],dout6[2],sp6[4],dout6[3],sout6[3],sp6[3]);
divide_module m1641(1'b0,d[4],dout6[3],sp6[5],dout6[4],sout6[4],sp6[4]);
divide_module m1651(1'b0,d[5],dout6[4],sp6[6],dout6[5],sout6[5],sp6[5]);
divide_module m1661(1'b0,d[6],dout6[5],sp6[7],dout6[6],sout6[6],sp6[6]);
divide_module m1671(1'b0,d[7],dout6[6],sp6[8],dout6[7],sout6[7],sp6[7]);
divide_module m1681(1'b0,d[8],dout6[7],sp6[9],dout6[8],sout6[8],sp6[8]);
divide_module m1691(1'b0,d[9],dout6[8],sp6[10],dout6[9],sout6[9],sp6[9]);
divide_module m1701(1'b0,d[10],dout6[9],sp6[11],dout6[10],sout6[10],sp6[10]);
divide_module m1711(1'b0,d[11],dout6[10],sp6[12],dout6[11],sout6[11],sp6[11]);
divide_module m1721(1'b0,d[12],dout6[11],sp6[13],dout6[12],sout6[12],sp6[12]);
divide_module m1731(1'b0,d[13],dout6[12],sp6[14],dout6[13],sout6[13],sp6[13]);
divide_module m1741(1'b0,d[14],dout6[13],sp6[15],dout6[14],sout6[14],sp6[14]);
divide_module m1751(1'b0,d[15],dout6[14],sp6[16],dout6[15],sout6[15],sp6[15]);
divide_module m1761(1'b0,d[16],dout6[15],sp6[17],dout6[16],sout6[16],sp6[16]);
divide_module m1771(1'b0,d[17],dout6[16],sp6[18],dout6[17],sout6[17],sp6[17]);
divide_module m1781(1'b0,d[18],dout6[17],sp6[19],dout6[18],sout6[18],sp6[18]);
divide_module m1791(1'b0,d[19],dout6[18],sp6[20],dout6[19],sout6[19],sp6[19]);
divide_module m1801(1'b0,d[20],dout6[19],sp6[21],dout6[20],sout6[20],sp6[20]);
divide_module m1811(1'b0,d[21],dout6[20],sp6[22],dout6[21],sout6[21],sp6[21]);
divide_module m1821(1'b0,d[22],dout6[21],sp6[23],dout6[22],sout6[22],sp6[22]);
divide_module m1831(1'b0,d[23],dout6[22],sp6[24],dout6[23],sout6[23],sp6[23]);
divide_module m1841(1'b0,d[24],dout6[23],sp6[25],dout6[24],sout6[24],sp6[24]);
divide_module m1851(1'b0,d[25],dout6[24],sp6[26],dout6[25],sout6[25],sp6[25]);
divide_module m1861(1'b0,d[26],dout6[25],sp6[27],dout6[26],sout6[26],sp6[26]);
divide_module m1871(1'b0,d[27],dout6[26],sp6[28],dout6[27],sout6[27],sp6[27]);
divide_module m1881(1'b0,d[28],dout6[27],sp6[29],dout6[28],sout6[28],sp6[28]);
divide_module m1891(1'b0,d[29],dout6[28],sp6[30],dout6[29],sout6[29],sp6[29]);
divide_module m1901(1'b0,d[30],dout6[29],~dout6[30],dout6[30],sout6[30],sp6[30]);

divide_module m1602(D[23],d[0],1'b0,sp7[1],dout7[0],sout7[0],sp7[0]);
divide_module m1612(1'b0,d[1],dout7[0],sp7[2],dout7[1],sout7[1],sp7[1]);
divide_module m1622(1'b0,d[2],dout7[1],sp7[3],dout7[2],sout7[2],sp7[2]);
divide_module m1632(1'b0,d[3],dout7[2],sp7[4],dout7[3],sout7[3],sp7[3]);
divide_module m1642(1'b0,d[4],dout7[3],sp7[5],dout7[4],sout7[4],sp7[4]);
divide_module m1652(1'b0,d[5],dout7[4],sp7[6],dout7[5],sout7[5],sp7[5]);
divide_module m1662(1'b0,d[6],dout7[5],sp7[7],dout7[6],sout7[6],sp7[6]);
divide_module m1672(1'b0,d[7],dout7[6],sp7[8],dout7[7],sout7[7],sp7[7]);
divide_module m1682(1'b0,d[8],dout7[7],sp7[9],dout7[8],sout7[8],sp7[8]);
divide_module m1692(1'b0,d[9],dout7[8],sp7[10],dout7[9],sout7[9],sp7[9]);
divide_module m1702(1'b0,d[10],dout7[9],sp7[11],dout7[10],sout7[10],sp7[10]);
divide_module m1712(1'b0,d[11],dout7[10],sp7[12],dout7[11],sout7[11],sp7[11]);
divide_module m1722(1'b0,d[12],dout7[11],sp7[13],dout7[12],sout7[12],sp7[12]);
divide_module m1732(1'b0,d[13],dout7[12],sp7[14],dout7[13],sout7[13],sp7[13]);
divide_module m1742(1'b0,d[14],dout7[13],sp7[15],dout7[14],sout7[14],sp7[14]);
divide_module m1752(1'b0,d[15],dout7[14],sp7[16],dout7[15],sout7[15],sp7[15]);
divide_module m1762(1'b0,d[16],dout7[15],sp7[17],dout7[16],sout7[16],sp7[16]);
divide_module m1772(1'b0,d[17],dout7[16],sp7[18],dout7[17],sout7[17],sp7[17]);
divide_module m1782(1'b0,d[18],dout7[17],sp7[19],dout7[18],sout7[18],sp7[18]);
divide_module m1792(1'b0,d[19],dout7[18],sp7[20],dout7[19],sout7[19],sp7[19]);
divide_module m1802(1'b0,d[20],dout7[19],sp7[21],dout7[20],sout7[20],sp7[20]);
divide_module m1812(1'b0,d[21],dout7[20],sp7[22],dout7[21],sout7[21],sp7[21]);
divide_module m1822(1'b0,d[22],dout7[21],sp7[23],dout7[22],sout7[22],sp7[22]);
divide_module m1832(1'b0,d[23],dout7[22],sp7[24],dout7[23],sout7[23],sp7[23]);
divide_module m1842(1'b0,d[24],dout7[23],sp7[25],dout7[24],sout7[24],sp7[24]);
divide_module m1852(1'b0,d[25],dout7[24],sp7[26],dout7[25],sout7[25],sp7[25]);
divide_module m1862(1'b0,d[26],dout7[25],sp7[27],dout7[26],sout7[26],sp7[26]);
divide_module m1872(1'b0,d[27],dout7[26],sp7[28],dout7[27],sout7[27],sp7[27]);
divide_module m1882(1'b0,d[28],dout7[27],sp7[29],dout7[28],sout7[28],sp7[28]);
divide_module m1892(1'b0,d[29],dout7[28],sp7[30],dout7[29],sout7[29],sp7[29]);
divide_module m1902(1'b0,d[30],dout7[29],~dout7[30],dout7[30],sout7[30],sp7[30]);

divide_module m1603(D[22],d[0],1'b0,sp8[1],dout8[0],sout8[0],sp8[0]);
divide_module m1613(1'b0,d[1],dout8[0],sp8[2],dout8[1],sout8[1],sp8[1]);
divide_module m1623(1'b0,d[2],dout8[1],sp8[3],dout8[2],sout8[2],sp8[2]);
divide_module m1633(1'b0,d[3],dout8[2],sp8[4],dout8[3],sout8[3],sp8[3]);
divide_module m1643(1'b0,d[4],dout8[3],sp8[5],dout8[4],sout8[4],sp8[4]);
divide_module m1653(1'b0,d[5],dout8[4],sp8[6],dout8[5],sout8[5],sp8[5]);
divide_module m1663(1'b0,d[6],dout8[5],sp8[7],dout8[6],sout8[6],sp8[6]);
divide_module m1673(1'b0,d[7],dout8[6],sp8[8],dout8[7],sout8[7],sp8[7]);
divide_module m1683(1'b0,d[8],dout8[7],sp8[9],dout8[8],sout8[8],sp8[8]);
divide_module m1693(1'b0,d[9],dout8[8],sp8[10],dout8[9],sout8[9],sp8[9]);
divide_module m1703(1'b0,d[10],dout8[9],sp8[11],dout8[10],sout8[10],sp8[10]);
divide_module m1713(1'b0,d[11],dout8[10],sp8[12],dout8[11],sout8[11],sp8[11]);
divide_module m1723(1'b0,d[12],dout8[11],sp8[13],dout8[12],sout8[12],sp8[12]);
divide_module m1733(1'b0,d[13],dout8[12],sp8[14],dout8[13],sout8[13],sp8[13]);
divide_module m1743(1'b0,d[14],dout8[13],sp8[15],dout8[14],sout8[14],sp8[14]);
divide_module m1753(1'b0,d[15],dout8[14],sp8[16],dout8[15],sout8[15],sp8[15]);
divide_module m1763(1'b0,d[16],dout8[15],sp8[17],dout8[16],sout8[16],sp8[16]);
divide_module m1773(1'b0,d[17],dout8[16],sp8[18],dout8[17],sout8[17],sp8[17]);
divide_module m1783(1'b0,d[18],dout8[17],sp8[19],dout8[18],sout8[18],sp8[18]);
divide_module m1793(1'b0,d[19],dout8[18],sp8[20],dout8[19],sout8[19],sp8[19]);
divide_module m1803(1'b0,d[20],dout8[19],sp8[21],dout8[20],sout8[20],sp8[20]);
divide_module m1813(1'b0,d[21],dout8[20],sp8[22],dout8[21],sout8[21],sp8[21]);
divide_module m1823(1'b0,d[22],dout8[21],sp8[23],dout8[22],sout8[22],sp8[22]);
divide_module m1833(1'b0,d[23],dout8[22],sp8[24],dout8[23],sout8[23],sp8[23]);
divide_module m1843(1'b0,d[24],dout8[23],sp8[25],dout8[24],sout8[24],sp8[24]);
divide_module m1853(1'b0,d[25],dout8[24],sp8[26],dout8[25],sout8[25],sp8[25]);
divide_module m1863(1'b0,d[26],dout8[25],sp8[27],dout8[26],sout8[26],sp8[26]);
divide_module m1873(1'b0,d[27],dout8[26],sp8[28],dout8[27],sout8[27],sp8[27]);
divide_module m1883(1'b0,d[28],dout8[27],sp8[29],dout8[28],sout8[28],sp8[28]);
divide_module m1893(1'b0,d[29],dout8[28],sp8[30],dout8[29],sout8[29],sp8[29]);
divide_module m1903(1'b0,d[30],dout8[29],~dout8[30],dout8[30],sout8[30],sp8[30]);


divide_module m1604(D[21],d[0],1'b0,sp9[1],dout9[0],sout9[0],sp9[0]);
divide_module m1614(1'b0,d[1],dout9[0],sp9[2],dout9[1],sout9[1],sp9[1]);
divide_module m1624(1'b0,d[2],dout9[1],sp9[3],dout9[2],sout9[2],sp9[2]);
divide_module m1634(1'b0,d[3],dout9[2],sp9[4],dout9[3],sout9[3],sp9[3]);
divide_module m1644(1'b0,d[4],dout9[3],sp9[5],dout9[4],sout9[4],sp9[4]);
divide_module m1654(1'b0,d[5],dout9[4],sp9[6],dout9[5],sout9[5],sp9[5]);
divide_module m1664(1'b0,d[6],dout9[5],sp9[7],dout9[6],sout9[6],sp9[6]);
divide_module m1674(1'b0,d[7],dout9[6],sp9[8],dout9[7],sout9[7],sp9[7]);
divide_module m1684(1'b0,d[8],dout9[7],sp9[9],dout9[8],sout9[8],sp9[8]);
divide_module m1694(1'b0,d[9],dout9[8],sp9[10],dout9[9],sout9[9],sp9[9]);
divide_module m1704(1'b0,d[10],dout9[9],sp9[11],dout9[10],sout9[10],sp9[10]);
divide_module m1714(1'b0,d[11],dout9[10],sp9[12],dout9[11],sout9[11],sp9[11]);
divide_module m1724(1'b0,d[12],dout9[11],sp9[13],dout9[12],sout9[12],sp9[12]);
divide_module m1734(1'b0,d[13],dout9[12],sp9[14],dout9[13],sout9[13],sp9[13]);
divide_module m1744(1'b0,d[14],dout9[13],sp9[15],dout9[14],sout9[14],sp9[14]);
divide_module m1754(1'b0,d[15],dout9[14],sp9[16],dout9[15],sout9[15],sp9[15]);
divide_module m1764(1'b0,d[16],dout9[15],sp9[17],dout9[16],sout9[16],sp9[16]);
divide_module m1774(1'b0,d[17],dout9[16],sp9[18],dout9[17],sout9[17],sp9[17]);
divide_module m1784(1'b0,d[18],dout9[17],sp9[19],dout9[18],sout9[18],sp9[18]);
divide_module m1794(1'b0,d[19],dout9[18],sp9[20],dout9[19],sout9[19],sp9[19]);
divide_module m1804(1'b0,d[20],dout9[19],sp9[21],dout9[20],sout9[20],sp9[20]);
divide_module m1814(1'b0,d[21],dout9[20],sp9[22],dout9[21],sout9[21],sp9[21]);
divide_module m1824(1'b0,d[22],dout9[21],sp9[23],dout9[22],sout9[22],sp9[22]);
divide_module m1834(1'b0,d[23],dout9[22],sp9[24],dout9[23],sout9[23],sp9[23]);
divide_module m1844(1'b0,d[24],dout9[23],sp9[25],dout9[24],sout9[24],sp9[24]);
divide_module m1854(1'b0,d[25],dout9[24],sp9[26],dout9[25],sout9[25],sp9[25]);
divide_module m1864(1'b0,d[26],dout9[25],sp9[27],dout9[26],sout9[26],sp9[26]);
divide_module m1874(1'b0,d[27],dout9[26],sp9[28],dout9[27],sout9[27],sp9[27]);
divide_module m1884(1'b0,d[28],dout9[27],sp9[29],dout9[28],sout9[28],sp9[28]);
divide_module m1894(1'b0,d[29],dout9[28],sp9[30],dout9[29],sout9[29],sp9[29]);
divide_module m1904(1'b0,d[30],dout9[29],~dout9[30],dout9[30],sout9[30],sp9[30]);

divide_module m1605(D[20],d[0],1'b0,sp10[1],dout10[0],sout10[0],sp10[0]);
divide_module m1615(1'b0,d[1],dout10[0],sp10[2],dout10[1],sout10[1],sp10[1]);
divide_module m1625(1'b0,d[2],dout10[1],sp10[3],dout10[2],sout10[2],sp10[2]);
divide_module m1635(1'b0,d[3],dout10[2],sp10[4],dout10[3],sout10[3],sp10[3]);
divide_module m1645(1'b0,d[4],dout10[3],sp10[5],dout10[4],sout10[4],sp10[4]);
divide_module m1655(1'b0,d[5],dout10[4],sp10[6],dout10[5],sout10[5],sp10[5]);
divide_module m1665(1'b0,d[6],dout10[5],sp10[7],dout10[6],sout10[6],sp10[6]);
divide_module m1675(1'b0,d[7],dout10[6],sp10[8],dout10[7],sout10[7],sp10[7]);
divide_module m1685(1'b0,d[8],dout10[7],sp10[9],dout10[8],sout10[8],sp10[8]);
divide_module m1695(1'b0,d[9],dout10[8],sp10[10],dout10[9],sout10[9],sp10[9]);
divide_module m1705(1'b0,d[10],dout10[9],sp10[11],dout10[10],sout10[10],sp10[10]);
divide_module m1715(1'b0,d[11],dout10[10],sp10[12],dout10[11],sout10[11],sp10[11]);
divide_module m1725(1'b0,d[12],dout10[11],sp10[13],dout10[12],sout10[12],sp10[12]);
divide_module m1735(1'b0,d[13],dout10[12],sp10[14],dout10[13],sout10[13],sp10[13]);
divide_module m1745(1'b0,d[14],dout10[13],sp10[15],dout10[14],sout10[14],sp10[14]);
divide_module m1755(1'b0,d[15],dout10[14],sp10[16],dout10[15],sout10[15],sp10[15]);
divide_module m1765(1'b0,d[16],dout10[15],sp10[17],dout10[16],sout10[16],sp10[16]);
divide_module m1775(1'b0,d[17],dout10[16],sp10[18],dout10[17],sout10[17],sp10[17]);
divide_module m1785(1'b0,d[18],dout10[17],sp10[19],dout10[18],sout10[18],sp10[18]); 
divide_module m1795(1'b0,d[19],dout10[18],sp10[20],dout10[19],sout10[19],sp10[19]);
divide_module m1805(1'b0,d[20],dout10[19],sp10[21],dout10[20],sout10[20],sp10[20]);
divide_module m1815(1'b0,d[21],dout10[20],sp10[22],dout10[21],sout10[21],sp10[21]);
divide_module m1825(1'b0,d[22],dout10[21],sp10[23],dout10[22],sout10[22],sp10[22]);
divide_module m1835(1'b0,d[23],dout10[22],sp10[24],dout10[23],sout10[23],sp10[23]);
divide_module m1845(1'b0,d[24],dout10[23],sp10[25],dout10[24],sout10[24],sp10[24]);
divide_module m1855(1'b0,d[25],dout10[24],sp10[26],dout10[25],sout10[25],sp10[25]);
divide_module m1865(1'b0,d[26],dout10[25],sp10[27],dout10[26],sout10[26],sp10[26]);
divide_module m1875(1'b0,d[27],dout10[26],sp10[28],dout10[27],sout10[27],sp10[27]);
divide_module m1885(1'b0,d[28],dout10[27],sp10[29],dout10[28],sout10[28],sp10[28]);
divide_module m1895(1'b0,d[29],dout10[28],sp10[30],dout10[29],sout10[29],sp10[29]);
divide_module m1905(1'b0,d[30],dout10[29],~dout10[30],dout10[30],sout10[30],sp10[30]);

divide_module m1606(D[19],d[0],1'b0,sp11[1],dout11[0],sout11[0],sp11[0]);
divide_module m1616(1'b0,d[1],dout11[0],sp11[2],dout11[1],sout11[1],sp11[1]);
divide_module m1626(1'b0,d[2],dout11[1],sp11[3],dout11[2],sout11[2],sp11[2]);
divide_module m1636(1'b0,d[3],dout11[2],sp11[4],dout11[3],sout11[3],sp11[3]);
divide_module m1646(1'b0,d[4],dout11[3],sp11[5],dout11[4],sout11[4],sp11[4]);
divide_module m1656(1'b0,d[5],dout11[4],sp11[6],dout11[5],sout11[5],sp11[5]);
divide_module m1666(1'b0,d[6],dout11[5],sp11[7],dout11[6],sout11[6],sp11[6]);
divide_module m1676(1'b0,d[7],dout11[6],sp11[8],dout11[7],sout11[7],sp11[7]);
divide_module m1686(1'b0,d[8],dout11[7],sp11[9],dout11[8],sout11[8],sp11[8]);
divide_module m1696(1'b0,d[9],dout11[8],sp11[10],dout11[9],sout11[9],sp11[9]);
divide_module m1706(1'b0,d[10],dout11[9],sp11[11],dout11[10],sout11[10],sp11[10]);
divide_module m1716(1'b0,d[11],dout11[10],sp11[12],dout11[11],sout11[11],sp11[11]);
divide_module m1726(1'b0,d[12],dout11[11],sp11[13],dout11[12],sout11[12],sp11[12]);
divide_module m1736(1'b0,d[13],dout11[12],sp11[14],dout11[13],sout11[13],sp11[13]);
divide_module m1746(1'b0,d[14],dout11[13],sp11[15],dout11[14],sout11[14],sp11[14]);
divide_module m1756(1'b0,d[15],dout11[14],sp11[16],dout11[15],sout11[15],sp11[15]);
divide_module m1766(1'b0,d[16],dout11[15],sp11[17],dout11[16],sout11[16],sp11[16]);
divide_module m1776(1'b0,d[17],dout11[16],sp11[18],dout11[17],sout11[17],sp11[17]);
divide_module m1786(1'b0,d[18],dout11[17],sp11[19],dout11[18],sout11[18],sp11[18]);
divide_module m1796(1'b0,d[19],dout11[18],sp11[20],dout11[19],sout11[19],sp11[19]);
divide_module m1806(1'b0,d[20],dout11[19],sp11[21],dout11[20],sout11[20],sp11[20]);
divide_module m1816(1'b0,d[21],dout11[20],sp11[22],dout11[21],sout11[21],sp11[21]);
divide_module m1826(1'b0,d[22],dout11[21],sp11[23],dout11[22],sout11[22],sp11[22]);
divide_module m1836(1'b0,d[23],dout11[22],sp11[24],dout11[23],sout11[23],sp11[23]);
divide_module m1846(1'b0,d[24],dout11[23],sp11[25],dout11[24],sout11[24],sp11[24]);
divide_module m1856(1'b0,d[25],dout11[24],sp11[26],dout11[25],sout11[25],sp11[25]);
divide_module m1866(1'b0,d[26],dout11[25],sp11[27],dout11[26],sout11[26],sp11[26]);
divide_module m1876(1'b0,d[27],dout11[26],sp11[28],dout11[27],sout11[27],sp11[27]);
divide_module m1886(1'b0,d[28],dout11[27],sp11[29],dout11[28],sout11[28],sp11[28]);
divide_module m1896(1'b0,d[29],dout11[28],sp11[30],dout11[29],sout11[29],sp11[29]);
divide_module m1906(1'b0,d[30],dout11[29],~dout11[30],dout11[30],sout11[30],sp11[30]);

divide_module m1607(D[18],d[0],1'b0,sp12[1],dout12[0],sout12[0],sp12[0]);
divide_module m1617(1'b0,d[1],dout12[0],sp12[2],dout12[1],sout12[1],sp12[1]);
divide_module m1627(1'b0,d[2],dout12[1],sp12[3],dout12[2],sout12[2],sp12[2]);
divide_module m1637(1'b0,d[3],dout12[2],sp12[4],dout12[3],sout12[3],sp12[3]);
divide_module m1647(1'b0,d[4],dout12[3],sp12[5],dout12[4],sout12[4],sp12[4]);
divide_module m1657(1'b0,d[5],dout12[4],sp12[6],dout12[5],sout12[5],sp12[5]);
divide_module m1667(1'b0,d[6],dout12[5],sp12[7],dout12[6],sout12[6],sp12[6]);
divide_module m1677(1'b0,d[7],dout12[6],sp12[8],dout12[7],sout12[7],sp12[7]);
divide_module m1687(1'b0,d[8],dout12[7],sp12[9],dout12[8],sout12[8],sp12[8]);
divide_module m1697(1'b0,d[9],dout12[8],sp12[10],dout12[9],sout12[9],sp12[9]);
divide_module m1707(1'b0,d[10],dout12[9],sp12[11],dout12[10],sout12[10],sp12[10]);
divide_module m1717(1'b0,d[11],dout12[10],sp12[12],dout12[11],sout12[11],sp12[11]);
divide_module m1727(1'b0,d[12],dout12[11],sp12[13],dout12[12],sout12[12],sp12[12]);
divide_module m1737(1'b0,d[13],dout12[12],sp12[14],dout12[13],sout12[13],sp12[13]);
divide_module m1747(1'b0,d[14],dout12[13],sp12[15],dout12[14],sout12[14],sp12[14]);
divide_module m1757(1'b0,d[15],dout12[14],sp12[16],dout12[15],sout12[15],sp12[15]);
divide_module m1767(1'b0,d[16],dout12[15],sp12[17],dout12[16],sout12[16],sp12[16]);
divide_module m1777(1'b0,d[17],dout12[16],sp12[18],dout12[17],sout12[17],sp12[17]);
divide_module m1787(1'b0,d[18],dout12[17],sp12[19],dout12[18],sout12[18],sp12[18]);
divide_module m1797(1'b0,d[19],dout12[18],sp12[20],dout12[19],sout12[19],sp12[19]);
divide_module m1807(1'b0,d[20],dout12[19],sp12[21],dout12[20],sout12[20],sp12[20]);
divide_module m1817(1'b0,d[21],dout12[20],sp12[22],dout12[21],sout12[21],sp12[21]);
divide_module m1827(1'b0,d[22],dout12[21],sp12[23],dout12[22],sout12[22],sp12[22]);
divide_module m1837(1'b0,d[23],dout12[22],sp12[24],dout12[23],sout12[23],sp12[23]);
divide_module m1847(1'b0,d[24],dout12[23],sp12[25],dout12[24],sout12[24],sp12[24]);
divide_module m1857(1'b0,d[25],dout12[24],sp12[26],dout12[25],sout12[25],sp12[25]);
divide_module m1867(1'b0,d[26],dout12[25],sp12[27],dout12[26],sout12[26],sp12[26]);
divide_module m1877(1'b0,d[27],dout12[26],sp12[28],dout12[27],sout12[27],sp12[27]);
divide_module m1887(1'b0,d[28],dout12[27],sp12[29],dout12[28],sout12[28],sp12[28]);
divide_module m1897(1'b0,d[29],dout12[28],sp12[30],dout12[29],sout12[29],sp12[29]);
divide_module m1907(1'b0,d[30],dout12[29],~dout12[30],dout12[30],sout12[30],sp12[30]);

divide_module m1608(D[17],d[0],1'b0,sp13[1],dout13[0],sout13[0],sp13[0]);
divide_module m1618(1'b0,d[1],dout13[0],sp13[2],dout13[1],sout13[1],sp13[1]);
divide_module m1628(1'b0,d[2],dout13[1],sp13[3],dout13[2],sout13[2],sp13[2]);
divide_module m1638(1'b0,d[3],dout13[2],sp13[4],dout13[3],sout13[3],sp13[3]);
divide_module m1648(1'b0,d[4],dout13[3],sp13[5],dout13[4],sout13[4],sp13[4]);
divide_module m1658(1'b0,d[5],dout13[4],sp13[6],dout13[5],sout13[5],sp13[5]);
divide_module m1668(1'b0,d[6],dout13[5],sp13[7],dout13[6],sout13[6],sp13[6]);
divide_module m1678(1'b0,d[7],dout13[6],sp13[8],dout13[7],sout13[7],sp13[7]);
divide_module m1688(1'b0,d[8],dout13[7],sp13[9],dout13[8],sout13[8],sp13[8]);
divide_module m1698(1'b0,d[9],dout13[8],sp13[10],dout13[9],sout13[9],sp13[9]);
divide_module m1708(1'b0,d[10],dout13[9],sp13[11],dout13[10],sout13[10],sp13[10]);
divide_module m1718(1'b0,d[11],dout13[10],sp13[12],dout13[11],sout13[11],sp13[11]);
divide_module m1728(1'b0,d[12],dout13[11],sp13[13],dout13[12],sout13[12],sp13[12]);
divide_module m1738(1'b0,d[13],dout13[12],sp13[14],dout13[13],sout13[13],sp13[13]);
divide_module m1748(1'b0,d[14],dout13[13],sp13[15],dout13[14],sout13[14],sp13[14]);
divide_module m1758(1'b0,d[15],dout13[14],sp13[16],dout13[15],sout13[15],sp13[15]);
divide_module m1768(1'b0,d[16],dout13[15],sp13[17],dout13[16],sout13[16],sp13[16]);
divide_module m1778(1'b0,d[17],dout13[16],sp13[18],dout13[17],sout13[17],sp13[17]); 
divide_module m1788(1'b0,d[18],dout13[17],sp13[19],dout13[18],sout13[18],sp13[18]);
divide_module m1798(1'b0,d[19],dout13[18],sp13[20],dout13[19],sout13[19],sp13[19]);
divide_module m1808(1'b0,d[20],dout13[19],sp13[21],dout13[20],sout13[20],sp13[20]);
divide_module m1818(1'b0,d[21],dout13[20],sp13[22],dout13[21],sout13[21],sp13[21]);
divide_module m1828(1'b0,d[22],dout13[21],sp13[23],dout13[22],sout13[22],sp13[22]);
divide_module m1838(1'b0,d[23],dout13[22],sp13[24],dout13[23],sout13[23],sp13[23]);
divide_module m1848(1'b0,d[24],dout13[23],sp13[25],dout13[24],sout13[24],sp13[24]);
divide_module m1858(1'b0,d[25],dout13[24],sp13[26],dout13[25],sout13[25],sp13[25]);
divide_module m1868(1'b0,d[26],dout13[25],sp13[27],dout13[26],sout13[26],sp13[26]);
divide_module m1878(1'b0,d[27],dout13[26],sp13[28],dout13[27],sout13[27],sp13[27]);
divide_module m1888(1'b0,d[28],dout13[27],sp13[29],dout13[28],sout13[28],sp13[28]);
divide_module m1898(1'b0,d[29],dout13[28],sp13[30],dout13[29],sout13[29],sp13[29]);
divide_module m1908(1'b0,d[30],dout13[29],~dout13[30],dout13[30],sout13[30],sp13[30]);

divide_module m1609(D[16],d[0],1'b0,sp14[1],dout14[0],sout14[0],sp14[0]);
divide_module m1619(1'b0,d[1],dout14[0],sp14[2],dout14[1],sout14[1],sp14[1]);
divide_module m1629(1'b0,d[2],dout14[1],sp14[3],dout14[2],sout14[2],sp14[2]);
divide_module m1639(1'b0,d[3],dout14[2],sp14[4],dout14[3],sout14[3],sp14[3]);
divide_module m1649(1'b0,d[4],dout14[3],sp14[5],dout14[4],sout14[4],sp14[4]);
divide_module m1659(1'b0,d[5],dout14[4],sp14[6],dout14[5],sout14[5],sp14[5]);
divide_module m1669(1'b0,d[6],dout14[5],sp14[7],dout14[6],sout14[6],sp14[6]);
divide_module m1679(1'b0,d[7],dout14[6],sp14[8],dout14[7],sout14[7],sp14[7]);
divide_module m1689(1'b0,d[8],dout14[7],sp14[9],dout14[8],sout14[8],sp14[8]);
divide_module m1699(1'b0,d[9],dout14[8],sp14[10],dout14[9],sout14[9],sp14[9]);
divide_module m1709(1'b0,d[10],dout14[9],sp14[11],dout14[10],sout14[10],sp14[10]);
divide_module m1719(1'b0,d[11],dout14[10],sp14[12],dout14[11],sout14[11],sp14[11]);
divide_module m1729(1'b0,d[12],dout14[11],sp14[13],dout14[12],sout14[12],sp14[12]);
divide_module m1739(1'b0,d[13],dout14[12],sp14[14],dout14[13],sout14[13],sp14[13]);
divide_module m1749(1'b0,d[14],dout14[13],sp14[15],dout14[14],sout14[14],sp14[14]);
divide_module m1759(1'b0,d[15],dout14[14],sp14[16],dout14[15],sout14[15],sp14[15]);
divide_module m1769(1'b0,d[16],dout14[15],sp14[17],dout14[16],sout14[16],sp14[16]);
divide_module m1779(1'b0,d[17],dout14[16],sp14[18],dout14[17],sout14[17],sp14[17]);
divide_module m1789(1'b0,d[18],dout14[17],sp14[19],dout14[18],sout14[18],sp14[18]);
divide_module m1799(1'b0,d[19],dout14[18],sp14[20],dout14[19],sout14[19],sp14[19]);
divide_module m1809(1'b0,d[20],dout14[19],sp14[21],dout14[20],sout14[20],sp14[20]);
divide_module m1819(1'b0,d[21],dout14[20],sp14[22],dout14[21],sout14[21],sp14[21]);
divide_module m1829(1'b0,d[22],dout14[21],sp14[23],dout14[22],sout14[22],sp14[22]);
divide_module m1839(1'b0,d[23],dout14[22],sp14[24],dout14[23],sout14[23],sp14[23]);
divide_module m1849(1'b0,d[24],dout14[23],sp14[25],dout14[24],sout14[24],sp14[24]);
divide_module m1859(1'b0,d[25],dout14[24],sp14[26],dout14[25],sout14[25],sp14[25]);
divide_module m1869(1'b0,d[26],dout14[25],sp14[27],dout14[26],sout14[26],sp14[26]);
divide_module m1879(1'b0,d[27],dout14[26],sp14[28],dout14[27],sout14[27],sp14[27]);
divide_module m1889(1'b0,d[28],dout14[27],sp14[29],dout14[28],sout14[28],sp14[28]);
divide_module m1899(1'b0,d[29],dout14[28],sp14[30],dout14[29],sout14[29],sp14[29]);
divide_module m1909(1'b0,d[30],dout14[29],~dout14[30],dout14[30],sout14[30],sp14[30]);


divide_module m16010(D[15],d[0],1'b0,sp15[1],dout15[0],sout15[0],sp15[0]);
divide_module m16110(1'b0,d[1],dout15[0],sp15[2],dout15[1],sout15[1],sp15[1]);
divide_module m16210(1'b0,d[2],dout15[1],sp15[3],dout15[2],sout15[2],sp15[2]);
divide_module m16310(1'b0,d[3],dout15[2],sp15[4],dout15[3],sout15[3],sp15[3]);
divide_module m16410(1'b0,d[4],dout15[3],sp15[5],dout15[4],sout15[4],sp15[4]);
divide_module m16510(1'b0,d[5],dout15[4],sp15[6],dout15[5],sout15[5],sp15[5]);
divide_module m16610(1'b0,d[6],dout15[5],sp15[7],dout15[6],sout15[6],sp15[6]);
divide_module m16710(1'b0,d[7],dout15[6],sp15[8],dout15[7],sout15[7],sp15[7]);
divide_module m16810(1'b0,d[8],dout15[7],sp15[9],dout15[8],sout15[8],sp15[8]);
divide_module m16910(1'b0,d[9],dout15[8],sp15[10],dout15[9],sout15[9],sp15[9]);
divide_module m17010(1'b0,d[10],dout15[9],sp15[11],dout15[10],sout15[10],sp15[10]);
divide_module m17110(1'b0,d[11],dout15[10],sp15[12],dout15[11],sout15[11],sp15[11]);
divide_module m17210(1'b0,d[12],dout15[11],sp15[13],dout15[12],sout15[12],sp15[12]);
divide_module m17310(1'b0,d[13],dout15[12],sp15[14],dout15[13],sout15[13],sp15[13]);
divide_module m17410(1'b0,d[14],dout15[13],sp15[15],dout15[14],sout15[14],sp15[14]);
divide_module m17510(1'b0,d[15],dout15[14],sp15[16],dout15[15],sout15[15],sp15[15]);
divide_module m17610(1'b0,d[16],dout15[15],sp15[17],dout15[16],sout15[16],sp15[16]);
divide_module m17710(1'b0,d[17],dout15[16],sp15[18],dout15[17],sout15[17],sp15[17]);
divide_module m17810(1'b0,d[18],dout15[17],sp15[19],dout15[18],sout15[18],sp15[18]);
divide_module m17910(1'b0,d[19],dout15[18],sp15[20],dout15[19],sout15[19],sp15[19]);
divide_module m18010(1'b0,d[20],dout15[19],sp15[21],dout15[20],sout15[20],sp15[20]);
divide_module m18110(1'b0,d[21],dout15[20],sp15[22],dout15[21],sout15[21],sp15[21]);
divide_module m18210(1'b0,d[22],dout15[21],sp15[23],dout15[22],sout15[22],sp15[22]);
divide_module m18310(1'b0,d[23],dout15[22],sp15[24],dout15[23],sout15[23],sp15[23]);
divide_module m18410(1'b0,d[24],dout15[23],sp15[25],dout15[24],sout15[24],sp15[24]);
divide_module m18510(1'b0,d[25],dout15[24],sp15[26],dout15[25],sout15[25],sp15[25]);
divide_module m18610(1'b0,d[26],dout15[25],sp15[27],dout15[26],sout15[26],sp15[26]);
divide_module m18710(1'b0,d[27],dout15[26],sp15[28],dout15[27],sout15[27],sp15[27]);
divide_module m18810(1'b0,d[28],dout15[27],sp15[29],dout15[28],sout15[28],sp15[28]);
divide_module m18910(1'b0,d[29],dout15[28],sp15[30],dout15[29],sout15[29],sp15[29]);
divide_module m19010(1'b0,d[30],dout15[29],~dout15[30],dout15[30],sout15[30],sp15[30]);


divide_module m16011(D[14],d[0],1'b0,sp16[1],dout16[0],sout16[0],sp16[0]);
divide_module m16111(1'b0,d[1],dout16[0],sp16[2],dout16[1],sout16[1],sp16[1]);
divide_module m16211(1'b0,d[2],dout16[1],sp16[3],dout16[2],sout16[2],sp16[2]);
divide_module m16311(1'b0,d[3],dout16[2],sp16[4],dout16[3],sout16[3],sp16[3]);
divide_module m16411(1'b0,d[4],dout16[3],sp16[5],dout16[4],sout16[4],sp16[4]);
divide_module m16511(1'b0,d[5],dout16[4],sp16[6],dout16[5],sout16[5],sp16[5]);
divide_module m16611(1'b0,d[6],dout16[5],sp16[7],dout16[6],sout16[6],sp16[6]);
divide_module m16711(1'b0,d[7],dout16[6],sp16[8],dout16[7],sout16[7],sp16[7]);
divide_module m16811(1'b0,d[8],dout16[7],sp16[9],dout16[8],sout16[8],sp16[8]);
divide_module m16911(1'b0,d[9],dout16[8],sp16[10],dout16[9],sout16[9],sp16[9]);
divide_module m17011(1'b0,d[10],dout16[9],sp16[11],dout16[10],sout16[10],sp16[10]);
divide_module m17111(1'b0,d[11],dout16[10],sp16[12],dout16[11],sout16[11],sp16[11]);
divide_module m17211(1'b0,d[12],dout16[11],sp16[13],dout16[12],sout16[12],sp16[12]);
divide_module m17311(1'b0,d[13],dout16[12],sp16[14],dout16[13],sout16[13],sp16[13]);
divide_module m17411(1'b0,d[14],dout16[13],sp16[15],dout16[14],sout16[14],sp16[14]);
divide_module m17511(1'b0,d[15],dout16[14],sp16[16],dout16[15],sout16[15],sp16[15]);
divide_module m17611(1'b0,d[16],dout16[15],sp16[17],dout16[16],sout16[16],sp16[16]);
divide_module m17711(1'b0,d[17],dout16[16],sp16[18],dout16[17],sout16[17],sp16[17]);
divide_module m17811(1'b0,d[18],dout16[17],sp16[19],dout16[18],sout16[18],sp16[18]);
divide_module m17911(1'b0,d[19],dout16[18],sp16[20],dout16[19],sout16[19],sp16[19]);
divide_module m18011(1'b0,d[20],dout16[19],sp16[21],dout16[20],sout16[20],sp16[20]);
divide_module m18111(1'b0,d[21],dout16[20],sp16[22],dout16[21],sout16[21],sp16[21]);
divide_module m18211(1'b0,d[22],dout16[21],sp16[23],dout16[22],sout16[22],sp16[22]);
divide_module m18311(1'b0,d[23],dout16[22],sp16[24],dout16[23],sout16[23],sp16[23]);
divide_module m18411(1'b0,d[24],dout16[23],sp16[25],dout16[24],sout16[24],sp16[24]);
divide_module m18511(1'b0,d[25],dout16[24],sp16[26],dout16[25],sout16[25],sp16[25]);
divide_module m18611(1'b0,d[26],dout16[25],sp16[27],dout16[26],sout16[26],sp16[26]);
divide_module m18711(1'b0,d[27],dout16[26],sp16[28],dout16[27],sout16[27],sp16[27]);
divide_module m18811(1'b0,d[28],dout16[27],sp16[29],dout16[28],sout16[28],sp16[28]);
divide_module m18911(1'b0,d[29],dout16[28],sp16[30],dout16[29],sout16[29],sp16[29]);
divide_module m19011(1'b0,d[30],dout16[29],~dout16[30],dout16[30],sout16[30],sp16[30]);


divide_module m16012(D[13],d[0],1'b0,sp17[1],dout17[0],sout17[0],sp17[0]);
divide_module m16112(1'b0,d[1],dout17[0],sp17[2],dout17[1],sout17[1],sp17[1]);
divide_module m16212(1'b0,d[2],dout17[1],sp17[3],dout17[2],sout17[2],sp17[2]);
divide_module m16312(1'b0,d[3],dout17[2],sp17[4],dout17[3],sout17[3],sp17[3]);
divide_module m16412(1'b0,d[4],dout17[3],sp17[5],dout17[4],sout17[4],sp17[4]);
divide_module m16512(1'b0,d[5],dout17[4],sp17[6],dout17[5],sout17[5],sp17[5]);
divide_module m16612(1'b0,d[6],dout17[5],sp17[7],dout17[6],sout17[6],sp17[6]);
divide_module m16712(1'b0,d[7],dout17[6],sp17[8],dout17[7],sout17[7],sp17[7]);
divide_module m16812(1'b0,d[8],dout17[7],sp17[9],dout17[8],sout17[8],sp17[8]);
divide_module m16912(1'b0,d[9],dout17[8],sp17[10],dout17[9],sout17[9],sp17[9]);
divide_module m17012(1'b0,d[10],dout17[9],sp17[11],dout17[10],sout17[10],sp17[10]);
divide_module m17112(1'b0,d[11],dout17[10],sp17[12],dout17[11],sout17[11],sp17[11]);
divide_module m17212(1'b0,d[12],dout17[11],sp17[13],dout17[12],sout17[12],sp17[12]);
divide_module m17312(1'b0,d[13],dout17[12],sp17[14],dout17[13],sout17[13],sp17[13]);
divide_module m17412(1'b0,d[14],dout17[13],sp17[15],dout17[14],sout17[14],sp17[14]);
divide_module m17512(1'b0,d[15],dout17[14],sp17[16],dout17[15],sout17[15],sp17[15]);
divide_module m17612(1'b0,d[16],dout17[15],sp17[17],dout17[16],sout17[16],sp17[16]);
divide_module m17712(1'b0,d[17],dout17[16],sp17[18],dout17[17],sout17[17],sp17[17]);
divide_module m17812(1'b0,d[18],dout17[17],sp17[19],dout17[18],sout17[18],sp17[18]);
divide_module m17912(1'b0,d[19],dout17[18],sp17[20],dout17[19],sout17[19],sp17[19]);
divide_module m18012(1'b0,d[20],dout17[19],sp17[21],dout17[20],sout17[20],sp17[20]);
divide_module m18112(1'b0,d[21],dout17[20],sp17[22],dout17[21],sout17[21],sp17[21]);
divide_module m18212(1'b0,d[22],dout17[21],sp17[23],dout17[22],sout17[22],sp17[22]);
divide_module m18312(1'b0,d[23],dout17[22],sp17[24],dout17[23],sout17[23],sp17[23]);
divide_module m18412(1'b0,d[24],dout17[23],sp17[25],dout17[24],sout17[24],sp17[24]);
divide_module m18512(1'b0,d[25],dout17[24],sp17[26],dout17[25],sout17[25],sp17[25]);
divide_module m18612(1'b0,d[26],dout17[25],sp17[27],dout17[26],sout17[26],sp17[26]);
divide_module m18712(1'b0,d[27],dout17[26],sp17[28],dout17[27],sout17[27],sp17[27]);
divide_module m18812(1'b0,d[28],dout17[27],sp17[29],dout17[28],sout17[28],sp17[28]);
divide_module m18912(1'b0,d[29],dout17[28],sp17[30],dout17[29],sout17[29],sp17[29]);
divide_module m19012(1'b0,d[30],dout17[29],~dout17[30],dout17[30],sout17[30],sp17[30]);

divide_module m16013(D[12],d[0],1'b0,sp18[1],dout18[0],sout18[0],sp18[0]);
divide_module m16113(1'b0,d[1],dout18[0],sp18[2],dout18[1],sout18[1],sp18[1]);
divide_module m16213(1'b0,d[2],dout18[1],sp18[3],dout18[2],sout18[2],sp18[2]);
divide_module m16313(1'b0,d[3],dout18[2],sp18[4],dout18[3],sout18[3],sp18[3]);
divide_module m16413(1'b0,d[4],dout18[3],sp18[5],dout18[4],sout18[4],sp18[4]);
divide_module m16513(1'b0,d[5],dout18[4],sp18[6],dout18[5],sout18[5],sp18[5]);
divide_module m16613(1'b0,d[6],dout18[5],sp18[7],dout18[6],sout18[6],sp18[6]);
divide_module m16713(1'b0,d[7],dout18[6],sp18[8],dout18[7],sout18[7],sp18[7]);
divide_module m16813(1'b0,d[8],dout18[7],sp18[9],dout18[8],sout18[8],sp18[8]);
divide_module m16913(1'b0,d[9],dout18[8],sp18[10],dout18[9],sout18[9],sp18[9]);
divide_module m17013(1'b0,d[10],dout18[9],sp18[11],dout18[10],sout18[10],sp18[10]);
divide_module m17113(1'b0,d[11],dout18[10],sp18[12],dout18[11],sout18[11],sp18[11]);
divide_module m17213(1'b0,d[12],dout18[11],sp18[13],dout18[12],sout18[12],sp18[12]);
divide_module m17313(1'b0,d[13],dout18[12],sp18[14],dout18[13],sout18[13],sp18[13]);
divide_module m17413(1'b0,d[14],dout18[13],sp18[15],dout18[14],sout18[14],sp18[14]);
divide_module m17513(1'b0,d[15],dout18[14],sp18[16],dout18[15],sout18[15],sp18[15]);
divide_module m17613(1'b0,d[16],dout18[15],sp18[17],dout18[16],sout18[16],sp18[16]);
divide_module m17713(1'b0,d[17],dout18[16],sp18[18],dout18[17],sout18[17],sp18[17]);
divide_module m17813(1'b0,d[18],dout18[17],sp18[19],dout18[18],sout18[18],sp18[18]);
divide_module m17913(1'b0,d[19],dout18[18],sp18[20],dout18[19],sout18[19],sp18[19]);
divide_module m18013(1'b0,d[20],dout18[19],sp18[21],dout18[20],sout18[20],sp18[20]);
divide_module m18113(1'b0,d[21],dout18[20],sp18[22],dout18[21],sout18[21],sp18[21]);
divide_module m18213(1'b0,d[22],dout18[21],sp18[23],dout18[22],sout18[22],sp18[22]);
divide_module m18313(1'b0,d[23],dout18[22],sp18[24],dout18[23],sout18[23],sp18[23]);
divide_module m18413(1'b0,d[24],dout18[23],sp18[25],dout18[24],sout18[24],sp18[24]);
divide_module m18513(1'b0,d[25],dout18[24],sp18[26],dout18[25],sout18[25],sp18[25]);
divide_module m18613(1'b0,d[26],dout18[25],sp18[27],dout18[26],sout18[26],sp18[26]);
divide_module m18713(1'b0,d[27],dout18[26],sp18[28],dout18[27],sout18[27],sp18[27]);
divide_module m18813(1'b0,d[28],dout18[27],sp18[29],dout18[28],sout18[28],sp18[28]);
divide_module m18913(1'b0,d[29],dout18[28],sp18[30],dout18[29],sout18[29],sp18[29]);
divide_module m19013(1'b0,d[30],dout18[29],~dout18[30],dout18[30],sout18[30],sp18[30]);

divide_module m16014(D[11],d[0],1'b0,sp19[1],dout19[0],sout19[0],sp19[0]);
divide_module m16114(1'b0,d[1],dout19[0],sp19[2],dout19[1],sout19[1],sp19[1]);
divide_module m16214(1'b0,d[2],dout19[1],sp19[3],dout19[2],sout19[2],sp19[2]);
divide_module m16314(1'b0,d[3],dout19[2],sp19[4],dout19[3],sout19[3],sp19[3]);
divide_module m16414(1'b0,d[4],dout19[3],sp19[5],dout19[4],sout19[4],sp19[4]);
divide_module m16514(1'b0,d[5],dout19[4],sp19[6],dout19[5],sout19[5],sp19[5]);
divide_module m16614(1'b0,d[6],dout19[5],sp19[7],dout19[6],sout19[6],sp19[6]);
divide_module m16714(1'b0,d[7],dout19[6],sp19[8],dout19[7],sout19[7],sp19[7]);
divide_module m16814(1'b0,d[8],dout19[7],sp19[9],dout19[8],sout19[8],sp19[8]);
divide_module m16914(1'b0,d[9],dout19[8],sp19[10],dout19[9],sout19[9],sp19[9]);
divide_module m17014(1'b0,d[10],dout19[9],sp19[11],dout19[10],sout19[10],sp19[10]);
divide_module m17114(1'b0,d[11],dout19[10],sp19[12],dout19[11],sout19[11],sp19[11]);
divide_module m17214(1'b0,d[12],dout19[11],sp19[13],dout19[12],sout19[12],sp19[12]);
divide_module m17314(1'b0,d[13],dout19[12],sp19[14],dout19[13],sout19[13],sp19[13]);
divide_module m17414(1'b0,d[14],dout19[13],sp19[15],dout19[14],sout19[14],sp19[14]);
divide_module m17514(1'b0,d[15],dout19[14],sp19[16],dout19[15],sout19[15],sp19[15]);
divide_module m17614(1'b0,d[16],dout19[15],sp19[17],dout19[16],sout19[16],sp19[16]);
divide_module m17714(1'b0,d[17],dout19[16],sp19[18],dout19[17],sout19[17],sp19[17]);
divide_module m17814(1'b0,d[18],dout19[17],sp19[19],dout19[18],sout19[18],sp19[18]);
divide_module m17914(1'b0,d[19],dout19[18],sp19[20],dout19[19],sout19[19],sp19[19]);
divide_module m18014(1'b0,d[20],dout19[19],sp19[21],dout19[20],sout19[20],sp19[20]);
divide_module m18114(1'b0,d[21],dout19[20],sp19[22],dout19[21],sout19[21],sp19[21]);
divide_module m18214(1'b0,d[22],dout19[21],sp19[23],dout19[22],sout19[22],sp19[22]);
divide_module m18314(1'b0,d[23],dout19[22],sp19[24],dout19[23],sout19[23],sp19[23]);
divide_module m18414(1'b0,d[24],dout19[23],sp19[25],dout19[24],sout19[24],sp19[24]);
divide_module m18514(1'b0,d[25],dout19[24],sp19[26],dout19[25],sout19[25],sp19[25]);
divide_module m18614(1'b0,d[26],dout19[25],sp19[27],dout19[26],sout19[26],sp19[26]);
divide_module m18714(1'b0,d[27],dout19[26],sp19[28],dout19[27],sout19[27],sp19[27]);
divide_module m18814(1'b0,d[28],dout19[27],sp19[29],dout19[28],sout19[28],sp19[28]);
divide_module m18914(1'b0,d[29],dout19[28],sp19[30],dout19[29],sout19[29],sp19[29]);
divide_module m19014(1'b0,d[30],dout19[29],~dout19[30],dout19[30],sout19[30],sp19[30]);

divide_module m16015(D[10],d[0],1'b0,sp20[1],dout20[0],sout20[0],sp20[0]);
divide_module m16115(1'b0,d[1],dout20[0],sp20[2],dout20[1],sout20[1],sp20[1]);
divide_module m16215(1'b0,d[2],dout20[1],sp20[3],dout20[2],sout20[2],sp20[2]);
divide_module m16315(1'b0,d[3],dout20[2],sp20[4],dout20[3],sout20[3],sp20[3]);
divide_module m16415(1'b0,d[4],dout20[3],sp20[5],dout20[4],sout20[4],sp20[4]);
divide_module m16515(1'b0,d[5],dout20[4],sp20[6],dout20[5],sout20[5],sp20[5]);
divide_module m16615(1'b0,d[6],dout20[5],sp20[7],dout20[6],sout20[6],sp20[6]);
divide_module m16715(1'b0,d[7],dout20[6],sp20[8],dout20[7],sout20[7],sp20[7]);
divide_module m16815(1'b0,d[8],dout20[7],sp20[9],dout20[8],sout20[8],sp20[8]);
divide_module m16915(1'b0,d[9],dout20[8],sp20[10],dout20[9],sout20[9],sp20[9]);
divide_module m17015(1'b0,d[10],dout20[9],sp20[11],dout20[10],sout20[10],sp20[10]);
divide_module m17115(1'b0,d[11],dout20[10],sp20[12],dout20[11],sout20[11],sp20[11]);
divide_module m17215(1'b0,d[12],dout20[11],sp20[13],dout20[12],sout20[12],sp20[12]);
divide_module m17315(1'b0,d[13],dout20[12],sp20[14],dout20[13],sout20[13],sp20[13]);
divide_module m17415(1'b0,d[14],dout20[13],sp20[15],dout20[14],sout20[14],sp20[14]);
divide_module m17515(1'b0,d[15],dout20[14],sp20[16],dout20[15],sout20[15],sp20[15]);
divide_module m17615(1'b0,d[16],dout20[15],sp20[17],dout20[16],sout20[16],sp20[16]);
divide_module m17715(1'b0,d[17],dout20[16],sp20[18],dout20[17],sout20[17],sp20[17]);
divide_module m17815(1'b0,d[18],dout20[17],sp20[19],dout20[18],sout20[18],sp20[18]);
divide_module m17915(1'b0,d[19],dout20[18],sp20[20],dout20[19],sout20[19],sp20[19]);
divide_module m18015(1'b0,d[20],dout20[19],sp20[21],dout20[20],sout20[20],sp20[20]);
divide_module m18115(1'b0,d[21],dout20[20],sp20[22],dout20[21],sout20[21],sp20[21]);
divide_module m18215(1'b0,d[22],dout20[21],sp20[23],dout20[22],sout20[22],sp20[22]);
divide_module m18315(1'b0,d[23],dout20[22],sp20[24],dout20[23],sout20[23],sp20[23]);
divide_module m18415(1'b0,d[24],dout20[23],sp20[25],dout20[24],sout20[24],sp20[24]);
divide_module m18515(1'b0,d[25],dout20[24],sp20[26],dout20[25],sout20[25],sp20[25]);
divide_module m18615(1'b0,d[26],dout20[25],sp20[27],dout20[26],sout20[26],sp20[26]);
divide_module m18715(1'b0,d[27],dout20[26],sp20[28],dout20[27],sout20[27],sp20[27]);
divide_module m18815(1'b0,d[28],dout20[27],sp20[29],dout20[28],sout20[28],sp20[28]);
divide_module m18915(1'b0,d[29],dout20[28],sp20[30],dout20[29],sout20[29],sp20[29]);
divide_module m19015(1'b0,d[30],dout20[29],~dout20[30],dout20[30],sout20[30],sp20[30]);

divide_module m16016(D[9],d[0],1'b0,sp21[1],dout21[0],sout21[0],sp21[0]);
divide_module m16116(1'b0,d[1],dout21[0],sp21[2],dout21[1],sout21[1],sp21[1]);
divide_module m16216(1'b0,d[2],dout21[1],sp21[3],dout21[2],sout21[2],sp21[2]);
divide_module m16316(1'b0,d[3],dout21[2],sp21[4],dout21[3],sout21[3],sp21[3]);
divide_module m16416(1'b0,d[4],dout21[3],sp21[5],dout21[4],sout21[4],sp21[4]);
divide_module m16516(1'b0,d[5],dout21[4],sp21[6],dout21[5],sout21[5],sp21[5]);
divide_module m16616(1'b0,d[6],dout21[5],sp21[7],dout21[6],sout21[6],sp21[6]);
divide_module m16716(1'b0,d[7],dout21[6],sp21[8],dout21[7],sout21[7],sp21[7]);
divide_module m16816(1'b0,d[8],dout21[7],sp21[9],dout21[8],sout21[8],sp21[8]);
divide_module m16916(1'b0,d[9],dout21[8],sp21[10],dout21[9],sout21[9],sp21[9]);
divide_module m17016(1'b0,d[10],dout21[9],sp21[11],dout21[10],sout21[10],sp21[10]);
divide_module m17116(1'b0,d[11],dout21[10],sp21[12],dout21[11],sout21[11],sp21[11]);
divide_module m17216(1'b0,d[12],dout21[11],sp21[13],dout21[12],sout21[12],sp21[12]);
divide_module m17316(1'b0,d[13],dout21[12],sp21[14],dout21[13],sout21[13],sp21[13]);
divide_module m17416(1'b0,d[14],dout21[13],sp21[15],dout21[14],sout21[14],sp21[14]);
divide_module m17516(1'b0,d[15],dout21[14],sp21[16],dout21[15],sout21[15],sp21[15]);
divide_module m17616(1'b0,d[16],dout21[15],sp21[17],dout21[16],sout21[16],sp21[16]);
divide_module m17716(1'b0,d[17],dout21[16],sp21[18],dout21[17],sout21[17],sp21[17]);
divide_module m17816(1'b0,d[18],dout21[17],sp21[19],dout21[18],sout21[18],sp21[18]);
divide_module m17916(1'b0,d[19],dout21[18],sp21[20],dout21[19],sout21[19],sp21[19]);
divide_module m18016(1'b0,d[20],dout21[19],sp21[21],dout21[20],sout21[20],sp21[20]);
divide_module m18116(1'b0,d[21],dout21[20],sp21[22],dout21[21],sout21[21],sp21[21]);
divide_module m18216(1'b0,d[22],dout21[21],sp21[23],dout21[22],sout21[22],sp21[22]);
divide_module m18316(1'b0,d[23],dout21[22],sp21[24],dout21[23],sout21[23],sp21[23]);
divide_module m18416(1'b0,d[24],dout21[23],sp21[25],dout21[24],sout21[24],sp21[24]);
divide_module m18516(1'b0,d[25],dout21[24],sp21[26],dout21[25],sout21[25],sp21[25]);
divide_module m18616(1'b0,d[26],dout21[25],sp21[27],dout21[26],sout21[26],sp21[26]);
divide_module m18716(1'b0,d[27],dout21[26],sp21[28],dout21[27],sout21[27],sp21[27]);
divide_module m18816(1'b0,d[28],dout21[27],sp21[29],dout21[28],sout21[28],sp21[28]);
divide_module m18916(1'b0,d[29],dout21[28],sp21[30],dout21[29],sout21[29],sp21[29]);
divide_module m19016(1'b0,d[30],dout21[29],~dout21[30],dout21[30],sout21[30],sp21[30]);

divide_module m16017(D[8],d[0],1'b0,sp22[1],dout22[0],sout22[0],sp22[0]);
divide_module m16117(1'b0,d[1],dout22[0],sp22[2],dout22[1],sout22[1],sp22[1]);
divide_module m16217(1'b0,d[2],dout22[1],sp22[3],dout22[2],sout22[2],sp22[2]);
divide_module m16317(1'b0,d[3],dout22[2],sp22[4],dout22[3],sout22[3],sp22[3]);
divide_module m16417(1'b0,d[4],dout22[3],sp22[5],dout22[4],sout22[4],sp22[4]);
divide_module m16517(1'b0,d[5],dout22[4],sp22[6],dout22[5],sout22[5],sp22[5]);
divide_module m16617(1'b0,d[6],dout22[5],sp22[7],dout22[6],sout22[6],sp22[6]);
divide_module m16717(1'b0,d[7],dout22[6],sp22[8],dout22[7],sout22[7],sp22[7]);
divide_module m16817(1'b0,d[8],dout22[7],sp22[9],dout22[8],sout22[8],sp22[8]);
divide_module m16917(1'b0,d[9],dout22[8],sp22[10],dout22[9],sout22[9],sp22[9]);
divide_module m17017(1'b0,d[10],dout22[9],sp22[11],dout22[10],sout22[10],sp22[10]);
divide_module m17117(1'b0,d[11],dout22[10],sp22[12],dout22[11],sout22[11],sp22[11]);
divide_module m17217(1'b0,d[12],dout22[11],sp22[13],dout22[12],sout22[12],sp22[12]);
divide_module m17317(1'b0,d[13],dout22[12],sp22[14],dout22[13],sout22[13],sp22[13]);
divide_module m17417(1'b0,d[14],dout22[13],sp22[15],dout22[14],sout22[14],sp22[14]);
divide_module m17517(1'b0,d[15],dout22[14],sp22[16],dout22[15],sout22[15],sp22[15]);
divide_module m17617(1'b0,d[16],dout22[15],sp22[17],dout22[16],sout22[16],sp22[16]);
divide_module m17717(1'b0,d[17],dout22[16],sp22[18],dout22[17],sout22[17],sp22[17]);
divide_module m17817(1'b0,d[18],dout22[17],sp22[19],dout22[18],sout22[18],sp22[18]);
divide_module m17917(1'b0,d[19],dout22[18],sp22[20],dout22[19],sout22[19],sp22[19]);
divide_module m18017(1'b0,d[20],dout22[19],sp22[21],dout22[20],sout22[20],sp22[20]);
divide_module m18117(1'b0,d[21],dout22[20],sp22[22],dout22[21],sout22[21],sp22[21]);
divide_module m18217(1'b0,d[22],dout22[21],sp22[23],dout22[22],sout22[22],sp22[22]);
divide_module m18317(1'b0,d[23],dout22[22],sp22[24],dout22[23],sout22[23],sp22[23]);
divide_module m18417(1'b0,d[24],dout22[23],sp22[25],dout22[24],sout22[24],sp22[24]);
divide_module m18517(1'b0,d[25],dout22[24],sp22[26],dout22[25],sout22[25],sp22[25]);
divide_module m18617(1'b0,d[26],dout22[25],sp22[27],dout22[26],sout22[26],sp22[26]);
divide_module m18717(1'b0,d[27],dout22[26],sp22[28],dout22[27],sout22[27],sp22[27]);
divide_module m18817(1'b0,d[28],dout22[27],sp22[29],dout22[28],sout22[28],sp22[28]);
divide_module m18917(1'b0,d[29],dout22[28],sp22[30],dout22[29],sout22[29],sp22[29]);
divide_module m19017(1'b0,d[30],dout22[29],~dout22[30],dout22[30],sout22[30],sp22[30]);


divide_module m16018(D[7],d[0],1'b0,sp23[1],dout23[0],sout23[0],sp23[0]);
divide_module m16118(1'b0,d[1],dout23[0],sp23[2],dout23[1],sout23[1],sp23[1]);
divide_module m16218(1'b0,d[2],dout23[1],sp23[3],dout23[2],sout23[2],sp23[2]);
divide_module m16318(1'b0,d[3],dout23[2],sp23[4],dout23[3],sout23[3],sp23[3]);
divide_module m16418(1'b0,d[4],dout23[3],sp23[5],dout23[4],sout23[4],sp23[4]);
divide_module m16518(1'b0,d[5],dout23[4],sp23[6],dout23[5],sout23[5],sp23[5]);
divide_module m16618(1'b0,d[6],dout23[5],sp23[7],dout23[6],sout23[6],sp23[6]);
divide_module m16718(1'b0,d[7],dout23[6],sp23[8],dout23[7],sout23[7],sp23[7]);
divide_module m16818(1'b0,d[8],dout23[7],sp23[9],dout23[8],sout23[8],sp23[8]);
divide_module m16918(1'b0,d[9],dout23[8],sp23[10],dout23[9],sout23[9],sp23[9]);
divide_module m17018(1'b0,d[10],dout23[9],sp23[11],dout23[10],sout23[10],sp23[10]);
divide_module m17118(1'b0,d[11],dout23[10],sp23[12],dout23[11],sout23[11],sp23[11]);
divide_module m17218(1'b0,d[12],dout23[11],sp23[13],dout23[12],sout23[12],sp23[12]);
divide_module m17318(1'b0,d[13],dout23[12],sp23[14],dout23[13],sout23[13],sp23[13]);
divide_module m17418(1'b0,d[14],dout23[13],sp23[15],dout23[14],sout23[14],sp23[14]);
divide_module m17518(1'b0,d[15],dout23[14],sp23[16],dout23[15],sout23[15],sp23[15]);
divide_module m17618(1'b0,d[16],dout23[15],sp23[17],dout23[16],sout23[16],sp23[16]);
divide_module m17718(1'b0,d[17],dout23[16],sp23[18],dout23[17],sout23[17],sp23[17]);
divide_module m17818(1'b0,d[18],dout23[17],sp23[19],dout23[18],sout23[18],sp23[18]);
divide_module m17918(1'b0,d[19],dout23[18],sp23[20],dout23[19],sout23[19],sp23[19]);
divide_module m18018(1'b0,d[20],dout23[19],sp23[21],dout23[20],sout23[20],sp23[20]);
divide_module m18118(1'b0,d[21],dout23[20],sp23[22],dout23[21],sout23[21],sp23[21]);
divide_module m18218(1'b0,d[22],dout23[21],sp23[23],dout23[22],sout23[22],sp23[22]);
divide_module m18318(1'b0,d[23],dout23[22],sp23[24],dout23[23],sout23[23],sp23[23]);
divide_module m18418(1'b0,d[24],dout23[23],sp23[25],dout23[24],sout23[24],sp23[24]);
divide_module m18518(1'b0,d[25],dout23[24],sp23[26],dout23[25],sout23[25],sp23[25]);
divide_module m18618(1'b0,d[26],dout23[25],sp23[27],dout23[26],sout23[26],sp23[26]);
divide_module m18718(1'b0,d[27],dout23[26],sp23[28],dout23[27],sout23[27],sp23[27]);
divide_module m18818(1'b0,d[28],dout23[27],sp23[29],dout23[28],sout23[28],sp23[28]);
divide_module m18918(1'b0,d[29],dout23[28],sp23[30],dout23[29],sout23[29],sp23[29]);
divide_module m19018(1'b0,d[30],dout23[29],~dout23[30],dout23[30],sout23[30],sp23[30]);

divide_module m16019(D[6],d[0],1'b0,sp24[1],dout24[0],sout24[0],sp24[0]);
divide_module m16119(1'b0,d[1],dout24[0],sp24[2],dout24[1],sout24[1],sp24[1]);
divide_module m16219(1'b0,d[2],dout24[1],sp24[3],dout24[2],sout24[2],sp24[2]);
divide_module m16319(1'b0,d[3],dout24[2],sp24[4],dout24[3],sout24[3],sp24[3]);
divide_module m16419(1'b0,d[4],dout24[3],sp24[5],dout24[4],sout24[4],sp24[4]);
divide_module m16519(1'b0,d[5],dout24[4],sp24[6],dout24[5],sout24[5],sp24[5]);
divide_module m16619(1'b0,d[6],dout24[5],sp24[7],dout24[6],sout24[6],sp24[6]);
divide_module m16719(1'b0,d[7],dout24[6],sp24[8],dout24[7],sout24[7],sp24[7]);
divide_module m16819(1'b0,d[8],dout24[7],sp24[9],dout24[8],sout24[8],sp24[8]);
divide_module m16919(1'b0,d[9],dout24[8],sp24[10],dout24[9],sout24[9],sp24[9]);
divide_module m17019(1'b0,d[10],dout24[9],sp24[11],dout24[10],sout24[10],sp24[10]);
divide_module m17119(1'b0,d[11],dout24[10],sp24[12],dout24[11],sout24[11],sp24[11]);
divide_module m17219(1'b0,d[12],dout24[11],sp24[13],dout24[12],sout24[12],sp24[12]);
divide_module m17319(1'b0,d[13],dout24[12],sp24[14],dout24[13],sout24[13],sp24[13]);
divide_module m17419(1'b0,d[14],dout24[13],sp24[15],dout24[14],sout24[14],sp24[14]);
divide_module m17519(1'b0,d[15],dout24[14],sp24[16],dout24[15],sout24[15],sp24[15]);
divide_module m17619(1'b0,d[16],dout24[15],sp24[17],dout24[16],sout24[16],sp24[16]);
divide_module m17719(1'b0,d[17],dout24[16],sp24[18],dout24[17],sout24[17],sp24[17]);
divide_module m17819(1'b0,d[18],dout24[17],sp24[19],dout24[18],sout24[18],sp24[18]);
divide_module m17919(1'b0,d[19],dout24[18],sp24[20],dout24[19],sout24[19],sp24[19]);
divide_module m18019(1'b0,d[20],dout24[19],sp24[21],dout24[20],sout24[20],sp24[20]);
divide_module m18119(1'b0,d[21],dout24[20],sp24[22],dout24[21],sout24[21],sp24[21]);
divide_module m18219(1'b0,d[22],dout24[21],sp24[23],dout24[22],sout24[22],sp24[22]);
divide_module m18319(1'b0,d[23],dout24[22],sp24[24],dout24[23],sout24[23],sp24[23]);
divide_module m18419(1'b0,d[24],dout24[23],sp24[25],dout24[24],sout24[24],sp24[24]);
divide_module m18519(1'b0,d[25],dout24[24],sp24[26],dout24[25],sout24[25],sp24[25]);
divide_module m18619(1'b0,d[26],dout24[25],sp24[27],dout24[26],sout24[26],sp24[26]);
divide_module m18719(1'b0,d[27],dout24[26],sp24[28],dout24[27],sout24[27],sp24[27]);
divide_module m18819(1'b0,d[28],dout24[27],sp24[29],dout24[28],sout24[28],sp24[28]);
divide_module m18919(1'b0,d[29],dout24[28],sp24[30],dout24[29],sout24[29],sp24[29]);
divide_module m19019(1'b0,d[30],dout24[29],~dout24[30],dout24[30],sout24[30],sp24[30]);

divide_module m16020(D[5],d[0],1'b0,sp25[1],dout25[0],sout25[0],sp25[0]);
divide_module m16120(1'b0,d[1],dout25[0],sp25[2],dout25[1],sout25[1],sp25[1]);
divide_module m16220(1'b0,d[2],dout25[1],sp25[3],dout25[2],sout25[2],sp25[2]);
divide_module m16320(1'b0,d[3],dout25[2],sp25[4],dout25[3],sout25[3],sp25[3]);
divide_module m16420(1'b0,d[4],dout25[3],sp25[5],dout25[4],sout25[4],sp25[4]);
divide_module m16520(1'b0,d[5],dout25[4],sp25[6],dout25[5],sout25[5],sp25[5]);
divide_module m16620(1'b0,d[6],dout25[5],sp25[7],dout25[6],sout25[6],sp25[6]);
divide_module m16720(1'b0,d[7],dout25[6],sp25[8],dout25[7],sout25[7],sp25[7]);
divide_module m16820(1'b0,d[8],dout25[7],sp25[9],dout25[8],sout25[8],sp25[8]);
divide_module m16920(1'b0,d[9],dout25[8],sp25[10],dout25[9],sout25[9],sp25[9]);
divide_module m17020(1'b0,d[10],dout25[9],sp25[11],dout25[10],sout25[10],sp25[10]);
divide_module m17120(1'b0,d[11],dout25[10],sp25[12],dout25[11],sout25[11],sp25[11]);
divide_module m17220(1'b0,d[12],dout25[11],sp25[13],dout25[12],sout25[12],sp25[12]);
divide_module m17320(1'b0,d[13],dout25[12],sp25[14],dout25[13],sout25[13],sp25[13]);
divide_module m17420(1'b0,d[14],dout25[13],sp25[15],dout25[14],sout25[14],sp25[14]);
divide_module m17520(1'b0,d[15],dout25[14],sp25[16],dout25[15],sout25[15],sp25[15]);
divide_module m17620(1'b0,d[16],dout25[15],sp25[17],dout25[16],sout25[16],sp25[16]);
divide_module m17720(1'b0,d[17],dout25[16],sp25[18],dout25[17],sout25[17],sp25[17]);
divide_module m17820(1'b0,d[18],dout25[17],sp25[19],dout25[18],sout25[18],sp25[18]);
divide_module m17920(1'b0,d[19],dout25[18],sp25[20],dout25[19],sout25[19],sp25[19]);
divide_module m18020(1'b0,d[20],dout25[19],sp25[21],dout25[20],sout25[20],sp25[20]);
divide_module m18120(1'b0,d[21],dout25[20],sp25[22],dout25[21],sout25[21],sp25[21]);
divide_module m18220(1'b0,d[22],dout25[21],sp25[23],dout25[22],sout25[22],sp25[22]);
divide_module m18320(1'b0,d[23],dout25[22],sp25[24],dout25[23],sout25[23],sp25[23]);
divide_module m18420(1'b0,d[24],dout25[23],sp25[25],dout25[24],sout25[24],sp25[24]);
divide_module m18520(1'b0,d[25],dout25[24],sp25[26],dout25[25],sout25[25],sp25[25]);
divide_module m18620(1'b0,d[26],dout25[25],sp25[27],dout25[26],sout25[26],sp25[26]);
divide_module m18720(1'b0,d[27],dout25[26],sp25[28],dout25[27],sout25[27],sp25[27]);
divide_module m18820(1'b0,d[28],dout25[27],sp25[29],dout25[28],sout25[28],sp25[28]);
divide_module m18920(1'b0,d[29],dout25[28],sp25[30],dout25[29],sout25[29],sp25[29]);
divide_module m19020(1'b0,d[30],dout25[29],~dout25[30],dout25[30],sout25[30],sp25[30]);


divide_module m16021(D[4],d[0],1'b0,sp26[1],dout26[0],sout26[0],sp26[0]);
divide_module m16121(1'b0,d[1],dout26[0],sp26[2],dout26[1],sout26[1],sp26[1]);
divide_module m16221(1'b0,d[2],dout26[1],sp26[3],dout26[2],sout26[2],sp26[2]);
divide_module m16321(1'b0,d[3],dout26[2],sp26[4],dout26[3],sout26[3],sp26[3]);
divide_module m16421(1'b0,d[4],dout26[3],sp26[5],dout26[4],sout26[4],sp26[4]);
divide_module m16521(1'b0,d[5],dout26[4],sp26[6],dout26[5],sout26[5],sp26[5]);
divide_module m16621(1'b0,d[6],dout26[5],sp26[7],dout26[6],sout26[6],sp26[6]);
divide_module m16721(1'b0,d[7],dout26[6],sp26[8],dout26[7],sout26[7],sp26[7]);
divide_module m16821(1'b0,d[8],dout26[7],sp26[9],dout26[8],sout26[8],sp26[8]);
divide_module m16921(1'b0,d[9],dout26[8],sp26[10],dout26[9],sout26[9],sp26[9]);
divide_module m17021(1'b0,d[10],dout26[9],sp26[11],dout26[10],sout26[10],sp26[10]);
divide_module m17121(1'b0,d[11],dout26[10],sp26[12],dout26[11],sout26[11],sp26[11]);
divide_module m17221(1'b0,d[12],dout26[11],sp26[13],dout26[12],sout26[12],sp26[12]);
divide_module m17321(1'b0,d[13],dout26[12],sp26[14],dout26[13],sout26[13],sp26[13]);
divide_module m17421(1'b0,d[14],dout26[13],sp26[15],dout26[14],sout26[14],sp26[14]);
divide_module m17521(1'b0,d[15],dout26[14],sp26[16],dout26[15],sout26[15],sp26[15]);
divide_module m17621(1'b0,d[16],dout26[15],sp26[17],dout26[16],sout26[16],sp26[16]);
divide_module m17721(1'b0,d[17],dout26[16],sp26[18],dout26[17],sout26[17],sp26[17]);
divide_module m17821(1'b0,d[18],dout26[17],sp26[19],dout26[18],sout26[18],sp26[18]);
divide_module m17921(1'b0,d[19],dout26[18],sp26[20],dout26[19],sout26[19],sp26[19]);
divide_module m18021(1'b0,d[20],dout26[19],sp26[21],dout26[20],sout26[20],sp26[20]);
divide_module m18121(1'b0,d[21],dout26[20],sp26[22],dout26[21],sout26[21],sp26[21]);
divide_module m18221(1'b0,d[22],dout26[21],sp26[23],dout26[22],sout26[22],sp26[22]);
divide_module m18321(1'b0,d[23],dout26[22],sp26[24],dout26[23],sout26[23],sp26[23]);
divide_module m18421(1'b0,d[24],dout26[23],sp26[25],dout26[24],sout26[24],sp26[24]);
divide_module m18521(1'b0,d[25],dout26[24],sp26[26],dout26[25],sout26[25],sp26[25]);
divide_module m18621(1'b0,d[26],dout26[25],sp26[27],dout26[26],sout26[26],sp26[26]);
divide_module m18721(1'b0,d[27],dout26[26],sp26[28],dout26[27],sout26[27],sp26[27]);
divide_module m18821(1'b0,d[28],dout26[27],sp26[29],dout26[28],sout26[28],sp26[28]);
divide_module m18921(1'b0,d[29],dout26[28],sp26[30],dout26[29],sout26[29],sp26[29]);
divide_module m19021(1'b0,d[30],dout26[29],~dout26[30],dout26[30],sout26[30],sp26[30]);



divide_module m16022(D[3],d[0],1'b0,sp27[1],dout27[0],sout27[0],sp27[0]);
divide_module m16122(1'b0,d[1],dout27[0],sp27[2],dout27[1],sout27[1],sp27[1]);
divide_module m16222(1'b0,d[2],dout27[1],sp27[3],dout27[2],sout27[2],sp27[2]);
divide_module m16322(1'b0,d[3],dout27[2],sp27[4],dout27[3],sout27[3],sp27[3]);
divide_module m16422(1'b0,d[4],dout27[3],sp27[5],dout27[4],sout27[4],sp27[4]);
divide_module m16522(1'b0,d[5],dout27[4],sp27[6],dout27[5],sout27[5],sp27[5]);
divide_module m16622(1'b0,d[6],dout27[5],sp27[7],dout27[6],sout27[6],sp27[6]);
divide_module m16722(1'b0,d[7],dout27[6],sp27[8],dout27[7],sout27[7],sp27[7]);
divide_module m16822(1'b0,d[8],dout27[7],sp27[9],dout27[8],sout27[8],sp27[8]);
divide_module m16922(1'b0,d[9],dout27[8],sp27[10],dout27[9],sout27[9],sp27[9]);
divide_module m17022(1'b0,d[10],dout27[9],sp27[11],dout27[10],sout27[10],sp27[10]);
divide_module m17122(1'b0,d[11],dout27[10],sp27[12],dout27[11],sout27[11],sp27[11]);
divide_module m17222(1'b0,d[12],dout27[11],sp27[13],dout27[12],sout27[12],sp27[12]);
divide_module m17322(1'b0,d[13],dout27[12],sp27[14],dout27[13],sout27[13],sp27[13]);
divide_module m17422(1'b0,d[14],dout27[13],sp27[15],dout27[14],sout27[14],sp27[14]);
divide_module m17522(1'b0,d[15],dout27[14],sp27[16],dout27[15],sout27[15],sp27[15]);
divide_module m17622(1'b0,d[16],dout27[15],sp27[17],dout27[16],sout27[16],sp27[16]);
divide_module m17722(1'b0,d[17],dout27[16],sp27[18],dout27[17],sout27[17],sp27[17]);
divide_module m17822(1'b0,d[18],dout27[17],sp27[19],dout27[18],sout27[18],sp27[18]);
divide_module m17922(1'b0,d[19],dout27[18],sp27[20],dout27[19],sout27[19],sp27[19]);
divide_module m18022(1'b0,d[20],dout27[19],sp27[21],dout27[20],sout27[20],sp27[20]);
divide_module m18122(1'b0,d[21],dout27[20],sp27[22],dout27[21],sout27[21],sp27[21]);
divide_module m18222(1'b0,d[22],dout27[21],sp27[23],dout27[22],sout27[22],sp27[22]);
divide_module m18322(1'b0,d[23],dout27[22],sp27[24],dout27[23],sout27[23],sp27[23]);
divide_module m18422(1'b0,d[24],dout27[23],sp27[25],dout27[24],sout27[24],sp27[24]);
divide_module m18522(1'b0,d[25],dout27[24],sp27[26],dout27[25],sout27[25],sp27[25]);
divide_module m18622(1'b0,d[26],dout27[25],sp27[27],dout27[26],sout27[26],sp27[26]);
divide_module m18722(1'b0,d[27],dout27[26],sp27[28],dout27[27],sout27[27],sp27[27]);
divide_module m18822(1'b0,d[28],dout27[27],sp27[29],dout27[28],sout27[28],sp27[28]);
divide_module m18922(1'b0,d[29],dout27[28],sp27[30],dout27[29],sout27[29],sp27[29]);
divide_module m19022(1'b0,d[30],dout27[29],~dout27[30],dout27[30],sout27[30],sp27[30]);


divide_module m16023(D[2],d[0],1'b0,sp28[1],dout28[0],sout28[0],sp28[0]);
divide_module m16123(1'b0,d[1],dout28[0],sp28[2],dout28[1],sout28[1],sp28[1]);
divide_module m16223(1'b0,d[2],dout28[1],sp28[3],dout28[2],sout28[2],sp28[2]);
divide_module m16323(1'b0,d[3],dout28[2],sp28[4],dout28[3],sout28[3],sp28[3]);
divide_module m16423(1'b0,d[4],dout28[3],sp28[5],dout28[4],sout28[4],sp28[4]);
divide_module m16523(1'b0,d[5],dout28[4],sp28[6],dout28[5],sout28[5],sp28[5]);
divide_module m16623(1'b0,d[6],dout28[5],sp28[7],dout28[6],sout28[6],sp28[6]);
divide_module m16723(1'b0,d[7],dout28[6],sp28[8],dout28[7],sout28[7],sp28[7]);
divide_module m16823(1'b0,d[8],dout28[7],sp28[9],dout28[8],sout28[8],sp28[8]);
divide_module m16923(1'b0,d[9],dout28[8],sp28[10],dout28[9],sout28[9],sp28[9]);
divide_module m17023(1'b0,d[10],dout28[9],sp28[11],dout28[10],sout28[10],sp28[10]);
divide_module m17123(1'b0,d[11],dout28[10],sp28[12],dout28[11],sout28[11],sp28[11]);
divide_module m17223(1'b0,d[12],dout28[11],sp28[13],dout28[12],sout28[12],sp28[12]);
divide_module m17323(1'b0,d[13],dout28[12],sp28[14],dout28[13],sout28[13],sp28[13]);
divide_module m17423(1'b0,d[14],dout28[13],sp28[15],dout28[14],sout28[14],sp28[14]);
divide_module m17523(1'b0,d[15],dout28[14],sp28[16],dout28[15],sout28[15],sp28[15]);
divide_module m17623(1'b0,d[16],dout28[15],sp28[17],dout28[16],sout28[16],sp28[16]);
divide_module m17723(1'b0,d[17],dout28[16],sp28[18],dout28[17],sout28[17],sp28[17]);
divide_module m17823(1'b0,d[18],dout28[17],sp28[19],dout28[18],sout28[18],sp28[18]);
divide_module m17923(1'b0,d[19],dout28[18],sp28[20],dout28[19],sout28[19],sp28[19]);
divide_module m18023(1'b0,d[20],dout28[19],sp28[21],dout28[20],sout28[20],sp28[20]);
divide_module m18123(1'b0,d[21],dout28[20],sp28[22],dout28[21],sout28[21],sp28[21]);
divide_module m18223(1'b0,d[22],dout28[21],sp28[23],dout28[22],sout28[22],sp28[22]);
divide_module m18323(1'b0,d[23],dout28[22],sp28[24],dout28[23],sout28[23],sp28[23]);
divide_module m18423(1'b0,d[24],dout28[23],sp28[25],dout28[24],sout28[24],sp28[24]);
divide_module m18523(1'b0,d[25],dout28[24],sp28[26],dout28[25],sout28[25],sp28[25]);
divide_module m18623(1'b0,d[26],dout28[25],sp28[27],dout28[26],sout28[26],sp28[26]);
divide_module m18723(1'b0,d[27],dout28[26],sp28[28],dout28[27],sout28[27],sp28[27]);
divide_module m18823(1'b0,d[28],dout28[27],sp28[29],dout28[28],sout28[28],sp28[28]);
divide_module m18923(1'b0,d[29],dout28[28],sp28[30],dout28[29],sout28[29],sp28[29]);
divide_module m19023(1'b0,d[30],dout28[29],~dout28[30],dout28[30],sout28[30],sp28[30]);

divide_module m16024(D[3],d[0],1'b0,sp29[1],dout29[0],sout29[0],sp29[0]);
divide_module m16124(1'b0,d[1],dout29[0],sp29[2],dout29[1],sout29[1],sp29[1]);
divide_module m16224(1'b0,d[2],dout29[1],sp29[3],dout29[2],sout29[2],sp29[2]);
divide_module m16324(1'b0,d[3],dout29[2],sp29[4],dout29[3],sout29[3],sp29[3]);
divide_module m16424(1'b0,d[4],dout29[3],sp29[5],dout29[4],sout29[4],sp29[4]);
divide_module m16524(1'b0,d[5],dout29[4],sp29[6],dout29[5],sout29[5],sp29[5]);
divide_module m16624(1'b0,d[6],dout29[5],sp29[7],dout29[6],sout29[6],sp29[6]);
divide_module m16724(1'b0,d[7],dout29[6],sp29[8],dout29[7],sout29[7],sp29[7]);
divide_module m16824(1'b0,d[8],dout29[7],sp29[9],dout29[8],sout29[8],sp29[8]);
divide_module m16924(1'b0,d[9],dout29[8],sp29[10],dout29[9],sout29[9],sp29[9]);
divide_module m17024(1'b0,d[10],dout29[9],sp29[11],dout29[10],sout29[10],sp29[10]);
divide_module m17124(1'b0,d[11],dout29[10],sp29[12],dout29[11],sout29[11],sp29[11]);
divide_module m17224(1'b0,d[12],dout29[11],sp29[13],dout29[12],sout29[12],sp29[12]);
divide_module m17324(1'b0,d[13],dout29[12],sp29[14],dout29[13],sout29[13],sp29[13]);
divide_module m17424(1'b0,d[14],dout29[13],sp29[15],dout29[14],sout29[14],sp29[14]);
divide_module m17524(1'b0,d[15],dout29[14],sp29[16],dout29[15],sout29[15],sp29[15]);
divide_module m17624(1'b0,d[16],dout29[15],sp29[17],dout29[16],sout29[16],sp29[16]);
divide_module m17724(1'b0,d[17],dout29[16],sp29[18],dout29[17],sout29[17],sp29[17]);
divide_module m17824(1'b0,d[18],dout29[17],sp29[19],dout29[18],sout29[18],sp29[18]);
divide_module m17924(1'b0,d[19],dout29[18],sp29[20],dout29[19],sout29[19],sp29[19]);
divide_module m18024(1'b0,d[20],dout29[19],sp29[21],dout29[20],sout29[20],sp29[20]);
divide_module m18124(1'b0,d[21],dout29[20],sp29[22],dout29[21],sout29[21],sp29[21]);
divide_module m18224(1'b0,d[22],dout29[21],sp29[23],dout29[22],sout29[22],sp29[22]);
divide_module m18324(1'b0,d[23],dout29[22],sp29[24],dout29[23],sout29[23],sp29[23]);
divide_module m18424(1'b0,d[24],dout29[23],sp29[25],dout29[24],sout29[24],sp29[24]);
divide_module m18524(1'b0,d[25],dout29[24],sp29[26],dout29[25],sout29[25],sp29[25]);
divide_module m18624(1'b0,d[26],dout29[25],sp29[27],dout29[26],sout29[26],sp29[26]);
divide_module m18724(1'b0,d[27],dout29[26],sp29[28],dout29[27],sout29[27],sp29[27]);
divide_module m18824(1'b0,d[28],dout29[27],sp29[29],dout29[28],sout29[28],sp29[28]);
divide_module m18924(1'b0,d[29],dout29[28],sp29[30],dout29[29],sout29[29],sp29[29]);
divide_module m19024(1'b0,d[30],dout29[29],~dout29[30],dout29[30],sout29[30],sp29[30]);

divide_module m16025(D[3],d[0],1'b0,sp30[1],dout30[0],sout30[0],sp30[0]);
divide_module m16125(1'b0,d[1],dout30[0],sp30[2],dout30[1],sout30[1],sp30[1]);
divide_module m16225(1'b0,d[2],dout30[1],sp30[3],dout30[2],sout30[2],sp30[2]);
divide_module m16325(1'b0,d[3],dout30[2],sp30[4],dout30[3],sout30[3],sp30[3]);
divide_module m16425(1'b0,d[4],dout30[3],sp30[5],dout30[4],sout30[4],sp30[4]);
divide_module m16525(1'b0,d[5],dout30[4],sp30[6],dout30[5],sout30[5],sp30[5]);
divide_module m16625(1'b0,d[6],dout30[5],sp30[7],dout30[6],sout30[6],sp30[6]);
divide_module m16725(1'b0,d[7],dout30[6],sp30[8],dout30[7],sout30[7],sp30[7]);
divide_module m16825(1'b0,d[8],dout30[7],sp30[9],dout30[8],sout30[8],sp30[8]);
divide_module m16925(1'b0,d[9],dout30[8],sp30[10],dout30[9],sout30[9],sp30[9]);
divide_module m17025(1'b0,d[10],dout30[9],sp30[11],dout30[10],sout30[10],sp30[10]);
divide_module m17125(1'b0,d[11],dout30[10],sp30[12],dout30[11],sout30[11],sp30[11]);
divide_module m17225(1'b0,d[12],dout30[11],sp30[13],dout30[12],sout30[12],sp30[12]);
divide_module m17325(1'b0,d[13],dout30[12],sp30[14],dout30[13],sout30[13],sp30[13]);
divide_module m17425(1'b0,d[14],dout30[13],sp30[15],dout30[14],sout30[14],sp30[14]);
divide_module m17525(1'b0,d[15],dout30[14],sp30[16],dout30[15],sout30[15],sp30[15]);
divide_module m17625(1'b0,d[16],dout30[15],sp30[17],dout30[16],sout30[16],sp30[16]);
divide_module m17725(1'b0,d[17],dout30[16],sp30[18],dout30[17],sout30[17],sp30[17]);
divide_module m17825(1'b0,d[18],dout30[17],sp30[19],dout30[18],sout30[18],sp30[18]);
divide_module m17925(1'b0,d[19],dout30[18],sp30[20],dout30[19],sout30[19],sp30[19]);
divide_module m18025(1'b0,d[20],dout30[19],sp30[21],dout30[20],sout30[20],sp30[20]);
divide_module m18125(1'b0,d[21],dout30[20],sp30[22],dout30[21],sout30[21],sp30[21]);
divide_module m18225(1'b0,d[22],dout30[21],sp30[23],dout30[22],sout30[22],sp30[22]);
divide_module m18325(1'b0,d[23],dout30[22],sp30[24],dout30[23],sout30[23],sp30[23]);
divide_module m18425(1'b0,d[24],dout30[23],sp30[25],dout30[24],sout30[24],sp30[24]);
divide_module m18525(1'b0,d[25],dout30[24],sp30[26],dout30[25],sout30[25],sp30[25]);
divide_module m18625(1'b0,d[26],dout30[25],sp30[27],dout30[26],sout30[26],sp30[26]);
divide_module m18725(1'b0,d[27],dout30[26],sp30[28],dout30[27],sout30[27],sp30[27]);
divide_module m18825(1'b0,d[28],dout30[27],sp30[29],dout30[28],sout30[28],sp30[28]);
divide_module m18925(1'b0,d[29],dout30[28],sp30[30],dout30[29],sout30[29],sp30[29]);
divide_module m19025(1'b0,d[30],dout30[29],~dout30[30],dout30[30],sout30[30],sp30[30]);




assign q[30]=~dout[30];
assign q[29]=~dout1[31];
assign q[28]=~dout2[31];
assign q[27]=~dout3[31];
assign q[26]=~dout4[31];
assign q[25]=~dout5[31];
assign q[24]=~dout6[31];
assign q[23]=~dout7[31];
assign q[22]=~dout8[31];
assign q[21]=~dout9[31];
assign q[20]=~dout10[31];
assign q[19]=~dout11[31];
assign q[18]=~dout12[31];
assign q[17]=~dout13[31];
assign q[16]=~dout14[31];
assign q[15]=~dout15[31];
assign q[14]=~dout16[31];
assign q[13]=~dout17[31];
assign q[12]=~dout18[31];
assign q[11]=~dout19[31];
assign q[10]=~dout20[31];
assign q[9]=~dout21[31];
assign q[8]=~dout22[31];
assign q[7]=~dout23[31];
assign q[6]=~dout24[31];
assign q[5]=~dout25[31];
assign q[4]=~dout26[31];
assign q[3]=~dout27[31];
assign q[2]=~dout28[31];
assign q[1]=~dout29[31];
assign q[0]=~dout30[31];


endmodule